
module mainfsm ( clk, reset, .Op({\Op<1> , \Op<0> }), .Funct({\Funct<5> , 
        \Funct<4> , \Funct<3> , \Funct<2> , \Funct<1> , \Funct<0> }), IRWrite, 
        AdrSrc, .ALUSrcA({\ALUSrcA<1> , \ALUSrcA<0> }), .ALUSrcB({\ALUSrcB<1> , 
        \ALUSrcB<0> }), .ResultSrc({\ResultSrc<1> , \ResultSrc<0> }), NextPC, 
        RegW, MemW, Branch, ALUOp );
  input clk, reset, \Op<1> , \Op<0> , \Funct<5> , \Funct<4> , \Funct<3> ,
         \Funct<2> , \Funct<1> , \Funct<0> ;
  output IRWrite, AdrSrc, \ALUSrcA<1> , \ALUSrcA<0> , \ALUSrcB<1> ,
         \ALUSrcB<0> , \ResultSrc<1> , \ResultSrc<0> , NextPC, RegW, MemW,
         Branch, ALUOp;
  wire   \state<2> , \state<1> , \nextstate<3> , \nextstate<2> ,
         \nextstate<1> , \nextstate<0> , n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n2, n3, n4, n5, n8, n19, n20, n21, n22, n23, n27, n28, n29,
         n30;

  DFFRHQXL \state_reg<2>  ( .D(\nextstate<2> ), .CK(clk), .RN(n30), .Q(
        \state<2> ) );
  DFFRXL \state_reg<3>  ( .D(\nextstate<3> ), .CK(clk), .RN(n30), .Q(n22), 
        .QN(n23) );
  DFFRHQXL \state_reg<1>  ( .D(\nextstate<1> ), .CK(clk), .RN(n30), .Q(
        \state<1> ) );
  DFFRX1 \state_reg<0>  ( .D(\nextstate<0> ), .CK(clk), .RN(n30), .Q(n20), 
        .QN(n21) );
  AOI21XL U3 ( .A0(n10), .A1(n11), .B0(n12), .Y(\nextstate<2> ) );
  INVX20 U4 ( .A(\state<2> ), .Y(n29) );
  OAI32X4 U5 ( .A0(n27), .A1(n2), .A2(n8), .B0(n22), .B1(n9), .Y(
        \nextstate<3> ) );
  BUFX20 U6 ( .A(n5), .Y(\ALUSrcA<1> ) );
  BUFX8 U7 ( .A(n23), .Y(n3) );
  DLY1X1 U8 ( .A(\ALUSrcA<1> ), .Y(Branch) );
  AOI31XL U9 ( .A0(n2), .A1(n29), .A2(n4), .B0(\ALUSrcA<1> ), .Y(n18) );
  NOR2X4 U10 ( .A(n3), .B(n2), .Y(n5) );
  INVX1 U11 ( .A(\ALUSrcB<1> ), .Y(n8) );
  OAI21X1 U12 ( .A0(n2), .A1(n9), .B0(n18), .Y(\ALUSrcB<0> ) );
  BUFX8 U13 ( .A(n21), .Y(n2) );
  NAND2X4 U14 ( .A(n29), .B(n3), .Y(n12) );
  CLKBUFX8 U15 ( .A(\state<1> ), .Y(n4) );
  INVX1 U16 ( .A(n29), .Y(n19) );
  NOR2X1 U17 ( .A(n8), .B(n20), .Y(NextPC) );
  INVX1 U18 ( .A(n8), .Y(\ALUSrcA<0> ) );
  NOR2X4 U19 ( .A(n12), .B(n4), .Y(\ALUSrcB<1> ) );
  AOI31XL U20 ( .A0(n4), .A1(n29), .A2(n20), .B0(MemW), .Y(n17) );
  OAI2BB1X1 U21 ( .A0N(n2), .A1N(\Funct<0> ), .B0(n4), .Y(n10) );
  NAND2BXL U22 ( .AN(\ALUSrcA<1> ), .B(n8), .Y(\ResultSrc<1> ) );
  NAND2XL U23 ( .A(n19), .B(n4), .Y(n9) );
  AOI21XL U24 ( .A0(n2), .A1(n22), .B0(\ResultSrc<0> ), .Y(n16) );
  OAI22XL U25 ( .A0(n20), .A1(n12), .B0(n8), .B1(n15), .Y(\nextstate<0> ) );
  INVXL U26 ( .A(\Op<1> ), .Y(n27) );
  INVXL U27 ( .A(\Op<0> ), .Y(n28) );
  NAND3XL U28 ( .A(n28), .B(n27), .C(n20), .Y(n11) );
  NOR3XL U29 ( .A(n2), .B(n4), .C(n29), .Y(MemW) );
  INVX1 U30 ( .A(n9), .Y(ALUOp) );
  NOR3X1 U31 ( .A(n20), .B(n4), .C(n29), .Y(\ResultSrc<0> ) );
  INVX1 U32 ( .A(n16), .Y(RegW) );
  OAI21XL U33 ( .A0(\Funct<5> ), .A1(\Op<1> ), .B0(n28), .Y(n15) );
  OAI21XL U34 ( .A0(n8), .A1(n13), .B0(n14), .Y(\nextstate<1> ) );
  OAI21XL U35 ( .A0(\Op<0> ), .A1(n27), .B0(n20), .Y(n13) );
  NAND4BXL U36 ( .AN(n12), .B(\Funct<0> ), .C(n4), .D(n2), .Y(n14) );
  INVX1 U37 ( .A(reset), .Y(n30) );
  INVX1 U38 ( .A(n17), .Y(AdrSrc) );
  BUFX3 U39 ( .A(NextPC), .Y(IRWrite) );
endmodule


module decode ( clk, reset, .Op({\Op<1> , \Op<0> }), .Funct({\Funct<5> , 
        \Funct<4> , \Funct<3> , \Funct<2> , \Funct<1> , \Funct<0> }), .Rd({
        \Rd<3> , \Rd<2> , \Rd<1> , \Rd<0> }), .FlagW({\FlagW<1> , \FlagW<0> }), 
        PCS, NextPC, RegW, MemW, IRWrite, AdrSrc, .ResultSrc({\ResultSrc<1> , 
        \ResultSrc<0> }), .ALUSrcA({\ALUSrcA<1> , \ALUSrcA<0> }), .ALUSrcB({
        \ALUSrcB<1> , \ALUSrcB<0> }), .ImmSrc({\ImmSrc<1> , \ImmSrc<0> }), 
    .RegSrc({\RegSrc<1> , \RegSrc<0> }), .ALUControl({\ALUControl<1> , 
        \ALUControl<0> }) );
  input clk, reset, \Op<1> , \Op<0> , \Funct<5> , \Funct<4> , \Funct<3> ,
         \Funct<2> , \Funct<1> , \Funct<0> , \Rd<3> , \Rd<2> , \Rd<1> ,
         \Rd<0> ;
  output \FlagW<1> , \FlagW<0> , PCS, NextPC, RegW, MemW, IRWrite, AdrSrc,
         \ResultSrc<1> , \ResultSrc<0> , \ALUSrcA<1> , \ALUSrcA<0> ,
         \ALUSrcB<1> , \ALUSrcB<0> , \ImmSrc<1> , \ImmSrc<0> , \RegSrc<1> ,
         \RegSrc<0> , \ALUControl<1> , \ALUControl<0> ;
  wire   n23, n24, n25, n26, n27, n28, Branch, ALUOp, n5, n6, n7, n8, n10, n12,
         n14, n16, n18, n20, n22;

  mainfsm fsm ( .clk(clk), .reset(reset), .Op({\Op<1> , \Op<0> }), .Funct({
        \Funct<5> , \Funct<4> , \Funct<3> , \Funct<2> , \Funct<1> , \Funct<0> }), .IRWrite(n23), .AdrSrc(n24), .ALUSrcA({n26, n27}), .ALUSrcB({n28, 
        \ALUSrcB<0> }), .ResultSrc({n25, \ResultSrc<0> }), .RegW(RegW), .MemW(
        MemW), .Branch(Branch), .ALUOp(ALUOp) );
  INVX8 U3 ( .A(n26), .Y(n16) );
  INVX1 U4 ( .A(n16), .Y(\ALUSrcA<1> ) );
  INVX1 U5 ( .A(n27), .Y(n14) );
  INVX1 U6 ( .A(n14), .Y(\ALUSrcA<0> ) );
  BUFX1 U7 ( .A(\Op<0> ), .Y(\RegSrc<1> ) );
  BUFX1 U8 ( .A(\Op<1> ), .Y(\RegSrc<0> ) );
  INVX1 U9 ( .A(n12), .Y(\ALUSrcB<1> ) );
  INVX1 U10 ( .A(n28), .Y(n12) );
  INVX1 U11 ( .A(n10), .Y(\ResultSrc<1> ) );
  INVX1 U12 ( .A(n25), .Y(n10) );
  INVX1 U13 ( .A(ALUOp), .Y(n22) );
  INVX1 U14 ( .A(n20), .Y(NextPC) );
  INVX1 U15 ( .A(n20), .Y(IRWrite) );
  INVX1 U16 ( .A(n23), .Y(n20) );
  INVX1 U17 ( .A(n7), .Y(\FlagW<1> ) );
  INVX1 U18 ( .A(n18), .Y(AdrSrc) );
  AOI31X1 U19 ( .A0(RegW), .A1(\Rd<3> ), .A2(n6), .B0(Branch), .Y(n5) );
  AND3X2 U20 ( .A(\Rd<1> ), .B(\Rd<0> ), .C(\Rd<2> ), .Y(n6) );
  NOR2X1 U21 ( .A(\Funct<3> ), .B(\Funct<2> ), .Y(n8) );
  AOI2BB1X1 U22 ( .A0N(\Funct<4> ), .A1N(n8), .B0(n22), .Y(\ALUControl<1> ) );
  INVX1 U23 ( .A(n5), .Y(PCS) );
  AOI2BB1X1 U24 ( .A0N(\Funct<4> ), .A1N(\Funct<2> ), .B0(n22), .Y(
        \ALUControl<0> ) );
  NOR3X1 U25 ( .A(n7), .B(\Funct<4> ), .C(n8), .Y(\FlagW<0> ) );
  NAND2X1 U26 ( .A(ALUOp), .B(\Funct<0> ), .Y(n7) );
  INVX1 U27 ( .A(n24), .Y(n18) );
  BUFX3 U28 ( .A(\Op<1> ), .Y(\ImmSrc<1> ) );
  BUFX3 U29 ( .A(\Op<0> ), .Y(\ImmSrc<0> ) );
endmodule


module flopenr_WIDTH2_0 ( clk, reset, en, .d({\d<1> , \d<0> }), .q({\q<1> , 
        \q<0> }) );
  input clk, reset, en, \d<1> , \d<0> ;
  output \q<1> , \q<0> ;
  wire   n1, n3, n2, n4, n5, n6;

  DFFRHQX1 \q_reg<0>  ( .D(n2), .CK(clk), .RN(n6), .Q(\q<0> ) );
  DFFRHQXL \q_reg<1>  ( .D(n4), .CK(clk), .RN(n6), .Q(\q<1> ) );
  INVX1 U2 ( .A(n3), .Y(n4) );
  INVX1 U3 ( .A(n1), .Y(n2) );
  AOI22X4 U4 ( .A0(en), .A1(\d<0> ), .B0(\q<0> ), .B1(n5), .Y(n1) );
  AOI22X1 U5 ( .A0(\d<1> ), .A1(en), .B0(\q<1> ), .B1(n5), .Y(n3) );
  INVX1 U6 ( .A(en), .Y(n5) );
  INVX1 U7 ( .A(reset), .Y(n6) );
endmodule


module flopenr_WIDTH2_1 ( clk, reset, en, .d({\d<1> , \d<0> }), .q({\q<1> , 
        \q<0> }) );
  input clk, reset, en, \d<1> , \d<0> ;
  output \q<1> , \q<0> ;
  wire   n2, n4, n5, n6, n7, n8;

  DFFRHQXL \q_reg<1>  ( .D(n2), .CK(clk), .RN(n6), .Q(\q<1> ) );
  DFFRHQXL \q_reg<0>  ( .D(n4), .CK(clk), .RN(n6), .Q(\q<0> ) );
  INVX8 U2 ( .A(n8), .Y(n4) );
  AOI22X4 U3 ( .A0(en), .A1(\d<0> ), .B0(\q<0> ), .B1(n5), .Y(n8) );
  INVX1 U4 ( .A(en), .Y(n5) );
  INVX1 U5 ( .A(n7), .Y(n2) );
  AOI22X1 U6 ( .A0(\d<1> ), .A1(en), .B0(\q<1> ), .B1(n5), .Y(n7) );
  INVX1 U7 ( .A(reset), .Y(n6) );
endmodule


module condcheck ( .Cond({\Cond<3> , \Cond<2> , \Cond<1> , \Cond<0> }), 
    .Flags({\Flags<3> , \Flags<2> , \Flags<1> , \Flags<0> }), CondEx );
  input \Cond<3> , \Cond<2> , \Cond<1> , \Cond<0> , \Flags<3> , \Flags<2> ,
         \Flags<1> , \Flags<0> ;
  output CondEx;
  wire   n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20,
         n1, n2, n3, n4;

  OAI21XL U2 ( .A0(n6), .A1(n2), .B0(n7), .Y(CondEx) );
  AOI222X1 U3 ( .A0(\Cond<0> ), .A1(n14), .B0(n15), .B1(n16), .C0(\Cond<1> ), 
        .C1(n17), .Y(n6) );
  AOI32X1 U4 ( .A0(\Cond<1> ), .A1(n8), .A2(\Cond<2> ), .B0(n9), .B1(n2), .Y(
        n7) );
  NOR2X1 U5 ( .A(\Flags<2> ), .B(\Cond<0> ), .Y(n15) );
  XNOR2X1 U6 ( .A(n1), .B(\Cond<0> ), .Y(n13) );
  XOR2X1 U7 ( .A(\Flags<2> ), .B(\Cond<0> ), .Y(n12) );
  OAI32X1 U8 ( .A0(n3), .A1(\Cond<1> ), .A2(n10), .B0(\Cond<2> ), .B1(n11), 
        .Y(n9) );
  XNOR2X1 U9 ( .A(\Flags<3> ), .B(\Cond<0> ), .Y(n10) );
  AOI22X1 U10 ( .A0(n12), .A1(n4), .B0(\Cond<1> ), .B1(n13), .Y(n11) );
  INVX1 U11 ( .A(\Cond<1> ), .Y(n4) );
  XOR2X1 U12 ( .A(\Flags<0> ), .B(\Flags<3> ), .Y(n18) );
  INVX1 U13 ( .A(\Cond<2> ), .Y(n3) );
  OAI21XL U14 ( .A0(\Cond<0> ), .A1(n18), .B0(n3), .Y(n17) );
  OAI21XL U15 ( .A0(\Cond<1> ), .A1(n19), .B0(n20), .Y(n14) );
  AOI21X1 U16 ( .A0(n3), .A1(n1), .B0(\Flags<2> ), .Y(n19) );
  OAI21XL U17 ( .A0(\Cond<1> ), .A1(\Cond<2> ), .B0(n18), .Y(n20) );
  INVX1 U18 ( .A(\Flags<1> ), .Y(n1) );
  XOR2X1 U19 ( .A(\Flags<0> ), .B(\Cond<0> ), .Y(n8) );
  OAI32X1 U20 ( .A0(n1), .A1(\Cond<2> ), .A2(\Cond<1> ), .B0(n3), .B1(n18), 
        .Y(n16) );
  INVX1 U21 ( .A(\Cond<3> ), .Y(n2) );
endmodule


module flopr_WIDTH1 ( clk, reset, .d(\d<0> ), .q(\q<0> ) );
  input clk, reset, \d<0> ;
  output \q<0> ;
  wire   n1;

  DFFRHQXL \q_reg<0>  ( .D(\d<0> ), .CK(clk), .RN(n1), .Q(\q<0> ) );
  INVXL U3 ( .A(reset), .Y(n1) );
endmodule


module condlogic ( clk, reset, .Cond({\Cond<3> , \Cond<2> , \Cond<1> , 
        \Cond<0> }), .ALUFlags({\ALUFlags<3> , \ALUFlags<2> , \ALUFlags<1> , 
        \ALUFlags<0> }), .FlagW({\FlagW<1> , \FlagW<0> }), PCS, NextPC, RegW, 
        MemW, PCWrite, RegWrite, MemWrite );
  input clk, reset, \Cond<3> , \Cond<2> , \Cond<1> , \Cond<0> , \ALUFlags<3> ,
         \ALUFlags<2> , \ALUFlags<1> , \ALUFlags<0> , \FlagW<1> , \FlagW<0> ,
         PCS, NextPC, RegW, MemW;
  output PCWrite, RegWrite, MemWrite;
  wire   \FlagWrite<1> , \FlagWrite<0> , \Flags<3> , \Flags<2> , \Flags<1> ,
         \Flags<0> , CondEx, CondExDelayed, n2;

  flopenr_WIDTH2_0 flagreg1 ( .clk(clk), .reset(reset), .en(\FlagWrite<1> ), 
        .d({\ALUFlags<3> , \ALUFlags<2> }), .q({\Flags<3> , \Flags<2> }) );
  flopenr_WIDTH2_1 flagreg0 ( .clk(clk), .reset(reset), .en(\FlagWrite<0> ), 
        .d({\ALUFlags<1> , \ALUFlags<0> }), .q({\Flags<1> , \Flags<0> }) );
  condcheck cc ( .Cond({\Cond<3> , \Cond<2> , \Cond<1> , \Cond<0> }), .Flags({
        \Flags<3> , \Flags<2> , \Flags<1> , \Flags<0> }), .CondEx(CondEx) );
  flopr_WIDTH1 condreg ( .clk(clk), .reset(reset), .d(CondEx), .q(
        CondExDelayed) );
  AND2X2 U1 ( .A(\FlagW<1> ), .B(CondEx), .Y(\FlagWrite<1> ) );
  INVX1 U2 ( .A(n2), .Y(PCWrite) );
  AOI21X1 U3 ( .A0(PCS), .A1(CondExDelayed), .B0(NextPC), .Y(n2) );
  AND2X2 U4 ( .A(\FlagW<0> ), .B(CondEx), .Y(\FlagWrite<0> ) );
  AND2X2 U5 ( .A(RegW), .B(CondExDelayed), .Y(RegWrite) );
  AND2X2 U6 ( .A(MemW), .B(CondExDelayed), .Y(MemWrite) );
endmodule


module controller ( clk, reset, .Instr({\Instr<31> , \Instr<30> , \Instr<29> , 
        \Instr<28> , \Instr<27> , \Instr<26> , \Instr<25> , \Instr<24> , 
        \Instr<23> , \Instr<22> , \Instr<21> , \Instr<20> , \Instr<19> , 
        \Instr<18> , \Instr<17> , \Instr<16> , \Instr<15> , \Instr<14> , 
        \Instr<13> , \Instr<12> }), .ALUFlags({\ALUFlags<3> , \ALUFlags<2> , 
        \ALUFlags<1> , \ALUFlags<0> }), PCWrite, MemWrite, RegWrite, IRWrite, 
        AdrSrc, .RegSrc({\RegSrc<1> , \RegSrc<0> }), .ALUSrcA({\ALUSrcA<1> , 
        \ALUSrcA<0> }), .ALUSrcB({\ALUSrcB<1> , \ALUSrcB<0> }), .ResultSrc({
        \ResultSrc<1> , \ResultSrc<0> }), .ImmSrc({\ImmSrc<1> , \ImmSrc<0> }), 
    .ALUControl({\ALUControl<1> , \ALUControl<0> }) );
  input clk, reset, \Instr<31> , \Instr<30> , \Instr<29> , \Instr<28> ,
         \Instr<27> , \Instr<26> , \Instr<25> , \Instr<24> , \Instr<23> ,
         \Instr<22> , \Instr<21> , \Instr<20> , \Instr<19> , \Instr<18> ,
         \Instr<17> , \Instr<16> , \Instr<15> , \Instr<14> , \Instr<13> ,
         \Instr<12> , \ALUFlags<3> , \ALUFlags<2> , \ALUFlags<1> ,
         \ALUFlags<0> ;
  output PCWrite, MemWrite, RegWrite, IRWrite, AdrSrc, \RegSrc<1> ,
         \RegSrc<0> , \ALUSrcA<1> , \ALUSrcA<0> , \ALUSrcB<1> , \ALUSrcB<0> ,
         \ResultSrc<1> , \ResultSrc<0> , \ImmSrc<1> , \ImmSrc<0> ,
         \ALUControl<1> , \ALUControl<0> ;
  wire   n17, n18, n19, n20, n21, n22, n23, \FlagW<1> , \FlagW<0> , PCS, RegW,
         MemW, n2, n4, n6, n9, n11, n13, n14, n16;
  wire   SYNOPSYS_UNCONNECTED__0;

  decode dec ( .clk(clk), .reset(reset), .Op({\Instr<27> , \Instr<26> }), 
        .Funct({\Instr<25> , \Instr<24> , \Instr<23> , \Instr<22> , 
        \Instr<21> , \Instr<20> }), .Rd({\Instr<15> , \Instr<14> , \Instr<13> , 
        \Instr<12> }), .FlagW({\FlagW<1> , \FlagW<0> }), .PCS(PCS), .RegW(RegW), .MemW(MemW), .IRWrite(n18), .AdrSrc(n19), .ResultSrc({n22, \ResultSrc<0> }), 
        .ALUSrcA({n20, SYNOPSYS_UNCONNECTED__0}), .ALUSrcB({n21, \ALUSrcB<0> }), .ImmSrc({\ImmSrc<1> , \ImmSrc<0> }), .RegSrc({\RegSrc<1> , \RegSrc<0> }), 
        .ALUControl({n23, \ALUControl<0> }) );
  condlogic cl ( .clk(clk), .reset(reset), .Cond({\Instr<31> , \Instr<30> , 
        \Instr<29> , \Instr<28> }), .ALUFlags({\ALUFlags<3> , \ALUFlags<2> , 
        \ALUFlags<1> , \ALUFlags<0> }), .FlagW({\FlagW<1> , \FlagW<0> }), 
        .PCS(PCS), .NextPC(n14), .RegW(RegW), .MemW(MemW), .PCWrite(n17), 
        .RegWrite(RegWrite), .MemWrite(MemWrite) );
  INVX4 U1 ( .A(n21), .Y(n6) );
  INVX8 U2 ( .A(n6), .Y(\ALUSrcB<1> ) );
  INVX1 U3 ( .A(n6), .Y(\ALUSrcA<0> ) );
  INVX1 U4 ( .A(n9), .Y(\ALUSrcA<1> ) );
  INVX1 U5 ( .A(n20), .Y(n9) );
  INVX1 U6 ( .A(n4), .Y(\ResultSrc<1> ) );
  INVX1 U7 ( .A(n22), .Y(n4) );
  INVX1 U8 ( .A(n13), .Y(IRWrite) );
  INVX1 U9 ( .A(n18), .Y(n13) );
  INVX1 U10 ( .A(n16), .Y(PCWrite) );
  INVX1 U11 ( .A(n17), .Y(n16) );
  INVX1 U12 ( .A(n2), .Y(\ALUControl<1> ) );
  INVX1 U13 ( .A(n23), .Y(n2) );
  INVX1 U14 ( .A(n11), .Y(AdrSrc) );
  INVX1 U15 ( .A(n19), .Y(n11) );
  INVX1 U16 ( .A(n13), .Y(n14) );
endmodule


module flopenr_WIDTH32_0 ( clk, reset, en, .d({\d<31> , \d<30> , \d<29> , 
        \d<28> , \d<27> , \d<26> , \d<25> , \d<24> , \d<23> , \d<22> , \d<21> , 
        \d<20> , \d<19> , \d<18> , \d<17> , \d<16> , \d<15> , \d<14> , \d<13> , 
        \d<12> , \d<11> , \d<10> , \d<9> , \d<8> , \d<7> , \d<6> , \d<5> , 
        \d<4> , \d<3> , \d<2> , \d<1> , \d<0> }), .q({\q<31> , \q<30> , 
        \q<29> , \q<28> , \q<27> , \q<26> , \q<25> , \q<24> , \q<23> , \q<22> , 
        \q<21> , \q<20> , \q<19> , \q<18> , \q<17> , \q<16> , \q<15> , \q<14> , 
        \q<13> , \q<12> , \q<11> , \q<10> , \q<9> , \q<8> , \q<7> , \q<6> , 
        \q<5> , \q<4> , \q<3> , \q<2> , \q<1> , \q<0> }) );
  input clk, reset, en, \d<31> , \d<30> , \d<29> , \d<28> , \d<27> , \d<26> ,
         \d<25> , \d<24> , \d<23> , \d<22> , \d<21> , \d<20> , \d<19> ,
         \d<18> , \d<17> , \d<16> , \d<15> , \d<14> , \d<13> , \d<12> ,
         \d<11> , \d<10> , \d<9> , \d<8> , \d<7> , \d<6> , \d<5> , \d<4> ,
         \d<3> , \d<2> , \d<1> , \d<0> ;
  output \q<31> , \q<30> , \q<29> , \q<28> , \q<27> , \q<26> , \q<25> ,
         \q<24> , \q<23> , \q<22> , \q<21> , \q<20> , \q<19> , \q<18> ,
         \q<17> , \q<16> , \q<15> , \q<14> , \q<13> , \q<12> , \q<11> ,
         \q<10> , \q<9> , \q<8> , \q<7> , \q<6> , \q<5> , \q<4> , \q<3> ,
         \q<2> , \q<1> , \q<0> ;
  wire   n1, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n2, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43,
         n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57,
         n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71,
         n72, n73, n74, n75, n76;

  DFFRHQX1 \q_reg<1>  ( .D(n74), .CK(clk), .RN(n76), .Q(\q<1> ) );
  DFFRHQX1 \q_reg<0>  ( .D(n75), .CK(clk), .RN(n76), .Q(\q<0> ) );
  DFFRHQXL \q_reg<3>  ( .D(n72), .CK(clk), .RN(n2), .Q(\q<3> ) );
  DFFRHQXL \q_reg<2>  ( .D(n73), .CK(clk), .RN(n34), .Q(\q<2> ) );
  DFFRHQXL \q_reg<31>  ( .D(n44), .CK(clk), .RN(n2), .Q(\q<31> ) );
  DFFRHQXL \q_reg<8>  ( .D(n67), .CK(clk), .RN(n34), .Q(\q<8> ) );
  DFFRHQXL \q_reg<9>  ( .D(n66), .CK(clk), .RN(n34), .Q(\q<9> ) );
  DFFRHQXL \q_reg<10>  ( .D(n65), .CK(clk), .RN(n34), .Q(\q<10> ) );
  DFFRHQXL \q_reg<30>  ( .D(n45), .CK(clk), .RN(n2), .Q(\q<30> ) );
  DFFRHQXL \q_reg<29>  ( .D(n46), .CK(clk), .RN(n2), .Q(\q<29> ) );
  DFFRHQXL \q_reg<28>  ( .D(n47), .CK(clk), .RN(n2), .Q(\q<28> ) );
  DFFRHQXL \q_reg<27>  ( .D(n48), .CK(clk), .RN(n2), .Q(\q<27> ) );
  DFFRHQXL \q_reg<26>  ( .D(n49), .CK(clk), .RN(n2), .Q(\q<26> ) );
  DFFRHQXL \q_reg<25>  ( .D(n50), .CK(clk), .RN(n2), .Q(\q<25> ) );
  DFFRHQXL \q_reg<24>  ( .D(n51), .CK(clk), .RN(n2), .Q(\q<24> ) );
  DFFRHQXL \q_reg<23>  ( .D(n52), .CK(clk), .RN(n2), .Q(\q<23> ) );
  DFFRHQXL \q_reg<22>  ( .D(n53), .CK(clk), .RN(n2), .Q(\q<22> ) );
  DFFRHQXL \q_reg<21>  ( .D(n54), .CK(clk), .RN(n2), .Q(\q<21> ) );
  DFFRHQXL \q_reg<20>  ( .D(n55), .CK(clk), .RN(n2), .Q(\q<20> ) );
  DFFRHQXL \q_reg<19>  ( .D(n56), .CK(clk), .RN(n34), .Q(\q<19> ) );
  DFFRHQXL \q_reg<18>  ( .D(n57), .CK(clk), .RN(n34), .Q(\q<18> ) );
  DFFRHQXL \q_reg<17>  ( .D(n58), .CK(clk), .RN(n34), .Q(\q<17> ) );
  DFFRHQXL \q_reg<16>  ( .D(n59), .CK(clk), .RN(n34), .Q(\q<16> ) );
  DFFRHQXL \q_reg<15>  ( .D(n60), .CK(clk), .RN(n34), .Q(\q<15> ) );
  DFFRHQXL \q_reg<14>  ( .D(n61), .CK(clk), .RN(n34), .Q(\q<14> ) );
  DFFRHQXL \q_reg<13>  ( .D(n62), .CK(clk), .RN(n34), .Q(\q<13> ) );
  DFFRHQXL \q_reg<12>  ( .D(n63), .CK(clk), .RN(n34), .Q(\q<12> ) );
  DFFRHQXL \q_reg<11>  ( .D(n64), .CK(clk), .RN(n34), .Q(\q<11> ) );
  DFFRHQXL \q_reg<7>  ( .D(n68), .CK(clk), .RN(n2), .Q(\q<7> ) );
  DFFRHQXL \q_reg<6>  ( .D(n69), .CK(clk), .RN(n34), .Q(\q<6> ) );
  DFFRHQXL \q_reg<5>  ( .D(n70), .CK(clk), .RN(n2), .Q(\q<5> ) );
  DFFRHQXL \q_reg<4>  ( .D(n71), .CK(clk), .RN(n34), .Q(\q<4> ) );
  AOI22XL U2 ( .A0(\d<30> ), .A1(n41), .B0(\q<30> ), .B1(n39), .Y(n32) );
  AOI22XL U3 ( .A0(\d<29> ), .A1(n36), .B0(\q<29> ), .B1(n37), .Y(n31) );
  AOI22XL U4 ( .A0(\d<28> ), .A1(n36), .B0(\q<28> ), .B1(n37), .Y(n30) );
  AOI22XL U5 ( .A0(\d<27> ), .A1(en), .B0(\q<27> ), .B1(n37), .Y(n29) );
  AOI22XL U6 ( .A0(\d<26> ), .A1(en), .B0(\q<26> ), .B1(n37), .Y(n28) );
  AOI22XL U7 ( .A0(\d<25> ), .A1(n36), .B0(\q<25> ), .B1(n38), .Y(n27) );
  AOI22XL U8 ( .A0(\d<24> ), .A1(n42), .B0(\q<24> ), .B1(n38), .Y(n26) );
  AOI22XL U9 ( .A0(\d<23> ), .A1(n36), .B0(\q<23> ), .B1(n38), .Y(n25) );
  AOI22XL U10 ( .A0(\d<22> ), .A1(en), .B0(\q<22> ), .B1(n37), .Y(n24) );
  AOI22XL U11 ( .A0(\d<21> ), .A1(n36), .B0(\q<21> ), .B1(n38), .Y(n23) );
  AOI22XL U12 ( .A0(\d<20> ), .A1(en), .B0(\q<20> ), .B1(n38), .Y(n22) );
  AOI22XL U13 ( .A0(\d<19> ), .A1(n36), .B0(\q<19> ), .B1(n38), .Y(n21) );
  AOI22XL U14 ( .A0(\d<18> ), .A1(n36), .B0(\q<18> ), .B1(n37), .Y(n20) );
  AOI22XL U15 ( .A0(\d<17> ), .A1(n36), .B0(\q<17> ), .B1(n38), .Y(n19) );
  AOI22XL U16 ( .A0(\d<16> ), .A1(n36), .B0(\q<16> ), .B1(n37), .Y(n18) );
  AOI22XL U17 ( .A0(\d<15> ), .A1(n36), .B0(\q<15> ), .B1(n39), .Y(n17) );
  AOI22XL U18 ( .A0(\d<14> ), .A1(n36), .B0(\q<14> ), .B1(n39), .Y(n16) );
  AOI22XL U19 ( .A0(\d<13> ), .A1(n36), .B0(\q<13> ), .B1(n39), .Y(n15) );
  AOI22XL U20 ( .A0(\d<12> ), .A1(n36), .B0(\q<12> ), .B1(n39), .Y(n14) );
  AOI22XL U21 ( .A0(\d<11> ), .A1(n36), .B0(\q<11> ), .B1(n39), .Y(n13) );
  AOI22XL U22 ( .A0(\d<10> ), .A1(n36), .B0(\q<10> ), .B1(n39), .Y(n12) );
  AOI22XL U23 ( .A0(\d<9> ), .A1(n36), .B0(\q<9> ), .B1(n40), .Y(n11) );
  AOI22XL U24 ( .A0(\d<8> ), .A1(n36), .B0(\q<8> ), .B1(n40), .Y(n10) );
  AOI22XL U25 ( .A0(\d<7> ), .A1(n36), .B0(\q<7> ), .B1(n43), .Y(n9) );
  AOI22XL U26 ( .A0(\d<6> ), .A1(n42), .B0(\q<6> ), .B1(n43), .Y(n8) );
  AOI22XL U27 ( .A0(\d<5> ), .A1(n41), .B0(\q<5> ), .B1(n40), .Y(n7) );
  AOI22XL U28 ( .A0(\d<4> ), .A1(n36), .B0(\q<4> ), .B1(n40), .Y(n6) );
  AOI22XL U29 ( .A0(\d<3> ), .A1(n36), .B0(\q<3> ), .B1(n40), .Y(n5) );
  AOI22XL U30 ( .A0(\d<2> ), .A1(n41), .B0(\q<2> ), .B1(n40), .Y(n4) );
  AOI22XL U31 ( .A0(\d<1> ), .A1(n41), .B0(\q<1> ), .B1(n43), .Y(n3) );
  AOI22XL U32 ( .A0(n36), .A1(\d<0> ), .B0(\q<0> ), .B1(n43), .Y(n1) );
  CLKINVX3 U33 ( .A(n43), .Y(n36) );
  INVX1 U34 ( .A(n41), .Y(n40) );
  INVX1 U35 ( .A(n41), .Y(n39) );
  INVX1 U36 ( .A(n42), .Y(n38) );
  INVX1 U37 ( .A(n42), .Y(n37) );
  INVX1 U38 ( .A(n43), .Y(n41) );
  INVX1 U39 ( .A(n43), .Y(n42) );
  INVX1 U40 ( .A(en), .Y(n43) );
  CLKINVX3 U41 ( .A(n35), .Y(n34) );
  CLKINVX3 U42 ( .A(n35), .Y(n2) );
  INVX1 U43 ( .A(n76), .Y(n35) );
  INVX1 U44 ( .A(n33), .Y(n44) );
  AOI22X1 U45 ( .A0(\d<31> ), .A1(en), .B0(\q<31> ), .B1(n40), .Y(n33) );
  INVX1 U46 ( .A(n28), .Y(n49) );
  INVX1 U47 ( .A(n29), .Y(n48) );
  INVX1 U48 ( .A(n30), .Y(n47) );
  INVX1 U49 ( .A(n31), .Y(n46) );
  INVX1 U50 ( .A(n32), .Y(n45) );
  INVX1 U51 ( .A(n23), .Y(n54) );
  INVX1 U52 ( .A(n24), .Y(n53) );
  INVX1 U53 ( .A(n25), .Y(n52) );
  INVX1 U54 ( .A(n26), .Y(n51) );
  INVX1 U55 ( .A(n27), .Y(n50) );
  INVX1 U56 ( .A(n18), .Y(n59) );
  INVX1 U57 ( .A(n19), .Y(n58) );
  INVX1 U58 ( .A(n20), .Y(n57) );
  INVX1 U59 ( .A(n21), .Y(n56) );
  INVX1 U60 ( .A(n22), .Y(n55) );
  INVX1 U61 ( .A(n13), .Y(n64) );
  INVX1 U62 ( .A(n14), .Y(n63) );
  INVX1 U63 ( .A(n15), .Y(n62) );
  INVX1 U64 ( .A(n16), .Y(n61) );
  INVX1 U65 ( .A(n17), .Y(n60) );
  INVX1 U66 ( .A(n10), .Y(n67) );
  INVX1 U67 ( .A(n11), .Y(n66) );
  INVX1 U68 ( .A(n12), .Y(n65) );
  INVX1 U69 ( .A(n8), .Y(n69) );
  INVX1 U70 ( .A(n9), .Y(n68) );
  INVX1 U71 ( .A(n3), .Y(n74) );
  INVX1 U72 ( .A(n4), .Y(n73) );
  INVX1 U73 ( .A(n5), .Y(n72) );
  INVX1 U74 ( .A(n6), .Y(n71) );
  INVX1 U75 ( .A(n7), .Y(n70) );
  INVX1 U76 ( .A(n1), .Y(n75) );
  INVXL U77 ( .A(reset), .Y(n76) );
endmodule


module flopenr_WIDTH32_1 ( clk, reset, en, .d({\d<31> , \d<30> , \d<29> , 
        \d<28> , \d<27> , \d<26> , \d<25> , \d<24> , \d<23> , \d<22> , \d<21> , 
        \d<20> , \d<19> , \d<18> , \d<17> , \d<16> , \d<15> , \d<14> , \d<13> , 
        \d<12> , \d<11> , \d<10> , \d<9> , \d<8> , \d<7> , \d<6> , \d<5> , 
        \d<4> , \d<3> , \d<2> , \d<1> , \d<0> }), .q({\q<31> , \q<30> , 
        \q<29> , \q<28> , \q<27> , \q<26> , \q<25> , \q<24> , \q<23> , \q<22> , 
        \q<21> , \q<20> , \q<19> , \q<18> , \q<17> , \q<16> , \q<15> , \q<14> , 
        \q<13> , \q<12> , \q<11> , \q<10> , \q<9> , \q<8> , \q<7> , \q<6> , 
        \q<5> , \q<4> , \q<3> , \q<2> , \q<1> , \q<0> }) );
  input clk, reset, en, \d<31> , \d<30> , \d<29> , \d<28> , \d<27> , \d<26> ,
         \d<25> , \d<24> , \d<23> , \d<22> , \d<21> , \d<20> , \d<19> ,
         \d<18> , \d<17> , \d<16> , \d<15> , \d<14> , \d<13> , \d<12> ,
         \d<11> , \d<10> , \d<9> , \d<8> , \d<7> , \d<6> , \d<5> , \d<4> ,
         \d<3> , \d<2> , \d<1> , \d<0> ;
  output \q<31> , \q<30> , \q<29> , \q<28> , \q<27> , \q<26> , \q<25> ,
         \q<24> , \q<23> , \q<22> , \q<21> , \q<20> , \q<19> , \q<18> ,
         \q<17> , \q<16> , \q<15> , \q<14> , \q<13> , \q<12> , \q<11> ,
         \q<10> , \q<9> , \q<8> , \q<7> , \q<6> , \q<5> , \q<4> , \q<3> ,
         \q<2> , \q<1> , \q<0> ;
  wire   n111, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74,
         n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88,
         n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101,
         n102, n103, n104, n105, n106, n107, n108, n109, n110;

  DFFRHQXL \q_reg<25>  ( .D(n52), .CK(clk), .RN(n34), .Q(\q<25> ) );
  DFFRHQXL \q_reg<31>  ( .D(n46), .CK(clk), .RN(n34), .Q(\q<31> ) );
  DFFRHQX2 \q_reg<30>  ( .D(n47), .CK(clk), .RN(n34), .Q(\q<30> ) );
  DFFRHQXL \q_reg<21>  ( .D(n56), .CK(clk), .RN(n34), .Q(\q<21> ) );
  DFFRHQXL \q_reg<23>  ( .D(n54), .CK(clk), .RN(n34), .Q(\q<23> ) );
  DFFRHQXL \q_reg<19>  ( .D(n58), .CK(clk), .RN(n35), .Q(\q<19> ) );
  DFFRHQXL \q_reg<18>  ( .D(n59), .CK(clk), .RN(n35), .Q(\q<18> ) );
  DFFRHQX1 \q_reg<22>  ( .D(n55), .CK(clk), .RN(n34), .Q(\q<22> ) );
  DFFRHQX1 \q_reg<24>  ( .D(n53), .CK(clk), .RN(n34), .Q(\q<24> ) );
  DFFRHQXL \q_reg<17>  ( .D(n60), .CK(clk), .RN(n35), .Q(\q<17> ) );
  DFFRHQXL \q_reg<16>  ( .D(n61), .CK(clk), .RN(n35), .Q(\q<16> ) );
  DFFRHQX2 \q_reg<14>  ( .D(n63), .CK(clk), .RN(n35), .Q(\q<14> ) );
  DFFRHQX2 \q_reg<15>  ( .D(n62), .CK(clk), .RN(n35), .Q(\q<15> ) );
  DFFRHQXL \q_reg<11>  ( .D(n66), .CK(clk), .RN(n35), .Q(\q<11> ) );
  DFFRHQXL \q_reg<10>  ( .D(n67), .CK(clk), .RN(n35), .Q(\q<10> ) );
  DFFRHQX2 \q_reg<12>  ( .D(n65), .CK(clk), .RN(n35), .Q(\q<12> ) );
  DFFRHQX2 \q_reg<13>  ( .D(n64), .CK(clk), .RN(n35), .Q(\q<13> ) );
  DFFRHQXL \q_reg<9>  ( .D(n68), .CK(clk), .RN(n35), .Q(\q<9> ) );
  DFFRHQXL \q_reg<8>  ( .D(n69), .CK(clk), .RN(n35), .Q(\q<8> ) );
  DFFRHQXL \q_reg<7>  ( .D(n70), .CK(clk), .RN(n34), .Q(\q<7> ) );
  DFFRHQXL \q_reg<6>  ( .D(n71), .CK(clk), .RN(n35), .Q(\q<6> ) );
  DFFRHQXL \q_reg<5>  ( .D(n72), .CK(clk), .RN(n34), .Q(\q<5> ) );
  DFFRHQXL \q_reg<4>  ( .D(n73), .CK(clk), .RN(n35), .Q(\q<4> ) );
  DFFRHQX1 \q_reg<3>  ( .D(n74), .CK(clk), .RN(n34), .Q(\q<3> ) );
  DFFRHQX1 \q_reg<2>  ( .D(n75), .CK(clk), .RN(n35), .Q(\q<2> ) );
  DFFRHQX1 \q_reg<1>  ( .D(n76), .CK(clk), .RN(n78), .Q(\q<1> ) );
  DFFRHQX1 \q_reg<0>  ( .D(n77), .CK(clk), .RN(n78), .Q(\q<0> ) );
  DFFRHQX1 \q_reg<20>  ( .D(n57), .CK(clk), .RN(n34), .Q(\q<20> ) );
  DFFRHQX1 \q_reg<26>  ( .D(n51), .CK(clk), .RN(n34), .Q(\q<26> ) );
  DFFRHQX2 \q_reg<29>  ( .D(n48), .CK(clk), .RN(n34), .Q(\q<29> ) );
  DFFRHQX2 \q_reg<28>  ( .D(n49), .CK(clk), .RN(n34), .Q(\q<28> ) );
  DFFRHQXL \q_reg<27>  ( .D(n50), .CK(clk), .RN(n34), .Q(n111) );
  BUFX3 U2 ( .A(n111), .Y(\q<27> ) );
  AOI22XL U3 ( .A0(\d<26> ), .A1(n38), .B0(\q<26> ), .B1(n39), .Y(n84) );
  AOI22XL U4 ( .A0(\d<27> ), .A1(n38), .B0(\q<27> ), .B1(n39), .Y(n83) );
  AOI22XL U5 ( .A0(\d<8> ), .A1(n38), .B0(\q<8> ), .B1(n37), .Y(n102) );
  AOI22XL U6 ( .A0(\d<4> ), .A1(en), .B0(\q<4> ), .B1(n41), .Y(n106) );
  AOI22XL U7 ( .A0(\d<5> ), .A1(en), .B0(\q<5> ), .B1(n42), .Y(n105) );
  AOI22XL U8 ( .A0(\d<6> ), .A1(en), .B0(\q<6> ), .B1(n42), .Y(n104) );
  AOI22XL U9 ( .A0(\d<7> ), .A1(n43), .B0(\q<7> ), .B1(n42), .Y(n103) );
  AOI22XL U10 ( .A0(n43), .A1(\d<0> ), .B0(\q<0> ), .B1(n39), .Y(n110) );
  AOI22XL U11 ( .A0(\d<1> ), .A1(n38), .B0(\q<1> ), .B1(n37), .Y(n109) );
  AOI22XL U12 ( .A0(\d<2> ), .A1(n38), .B0(\q<2> ), .B1(n37), .Y(n108) );
  AOI22XL U13 ( .A0(\d<3> ), .A1(n38), .B0(\q<3> ), .B1(n37), .Y(n107) );
  CLKINVX3 U14 ( .A(n45), .Y(n38) );
  INVX1 U15 ( .A(n44), .Y(n42) );
  INVX1 U16 ( .A(n44), .Y(n41) );
  INVX1 U17 ( .A(n44), .Y(n40) );
  INVX1 U18 ( .A(n44), .Y(n39) );
  INVX1 U19 ( .A(n37), .Y(n43) );
  INVX1 U20 ( .A(n45), .Y(n44) );
  INVX1 U21 ( .A(n43), .Y(n45) );
  INVX1 U22 ( .A(en), .Y(n37) );
  CLKINVX3 U23 ( .A(n36), .Y(n35) );
  CLKINVX3 U24 ( .A(n36), .Y(n34) );
  INVX1 U25 ( .A(n78), .Y(n36) );
  INVX1 U26 ( .A(n82), .Y(n49) );
  AOI22X1 U27 ( .A0(\d<28> ), .A1(n38), .B0(\q<28> ), .B1(n39), .Y(n82) );
  INVX1 U28 ( .A(n81), .Y(n48) );
  AOI22X1 U29 ( .A0(\d<29> ), .A1(n38), .B0(\q<29> ), .B1(n39), .Y(n81) );
  INVX1 U30 ( .A(n95), .Y(n62) );
  AOI22X1 U31 ( .A0(\d<15> ), .A1(n38), .B0(\q<15> ), .B1(n42), .Y(n95) );
  INVX1 U32 ( .A(n97), .Y(n64) );
  AOI22X1 U33 ( .A0(\d<13> ), .A1(n44), .B0(\q<13> ), .B1(n40), .Y(n97) );
  INVX1 U34 ( .A(n96), .Y(n63) );
  AOI22X1 U35 ( .A0(\d<14> ), .A1(en), .B0(\q<14> ), .B1(n42), .Y(n96) );
  INVX1 U36 ( .A(n98), .Y(n65) );
  AOI22X1 U37 ( .A0(\d<12> ), .A1(n38), .B0(\q<12> ), .B1(n41), .Y(n98) );
  INVX1 U38 ( .A(n80), .Y(n47) );
  AOI22X1 U39 ( .A0(\d<30> ), .A1(n38), .B0(\q<30> ), .B1(n39), .Y(n80) );
  INVX1 U40 ( .A(n84), .Y(n51) );
  INVX1 U41 ( .A(n83), .Y(n50) );
  INVX1 U42 ( .A(n90), .Y(n57) );
  AOI22X1 U43 ( .A0(\d<20> ), .A1(n38), .B0(\q<20> ), .B1(n40), .Y(n90) );
  INVX1 U44 ( .A(n110), .Y(n77) );
  INVX1 U45 ( .A(n102), .Y(n69) );
  INVX1 U46 ( .A(n101), .Y(n68) );
  AOI22X1 U47 ( .A0(\d<9> ), .A1(n43), .B0(\q<9> ), .B1(n41), .Y(n101) );
  INVX1 U48 ( .A(n100), .Y(n67) );
  AOI22X1 U49 ( .A0(\d<10> ), .A1(en), .B0(\q<10> ), .B1(n41), .Y(n100) );
  INVX1 U50 ( .A(n99), .Y(n66) );
  AOI22X1 U51 ( .A0(\d<11> ), .A1(en), .B0(\q<11> ), .B1(n42), .Y(n99) );
  INVX1 U52 ( .A(n94), .Y(n61) );
  AOI22X1 U53 ( .A0(\d<16> ), .A1(n38), .B0(\q<16> ), .B1(n41), .Y(n94) );
  INVX1 U54 ( .A(n93), .Y(n60) );
  AOI22X1 U55 ( .A0(\d<17> ), .A1(n43), .B0(\q<17> ), .B1(n41), .Y(n93) );
  INVX1 U56 ( .A(n92), .Y(n59) );
  AOI22X1 U57 ( .A0(\d<18> ), .A1(n44), .B0(\q<18> ), .B1(n41), .Y(n92) );
  INVX1 U58 ( .A(n91), .Y(n58) );
  AOI22X1 U59 ( .A0(\d<19> ), .A1(n43), .B0(\q<19> ), .B1(n42), .Y(n91) );
  INVX1 U60 ( .A(n89), .Y(n56) );
  AOI22X1 U61 ( .A0(\d<21> ), .A1(n38), .B0(\q<21> ), .B1(n40), .Y(n89) );
  INVX1 U62 ( .A(n88), .Y(n55) );
  AOI22X1 U63 ( .A0(\d<22> ), .A1(n38), .B0(\q<22> ), .B1(n40), .Y(n88) );
  INVX1 U64 ( .A(n87), .Y(n54) );
  AOI22X1 U65 ( .A0(\d<23> ), .A1(n38), .B0(\q<23> ), .B1(n40), .Y(n87) );
  INVX1 U66 ( .A(n86), .Y(n53) );
  AOI22X1 U67 ( .A0(\d<24> ), .A1(n38), .B0(\q<24> ), .B1(n40), .Y(n86) );
  INVX1 U68 ( .A(n85), .Y(n52) );
  AOI22X1 U69 ( .A0(\d<25> ), .A1(n38), .B0(\q<25> ), .B1(n40), .Y(n85) );
  INVX1 U70 ( .A(n79), .Y(n46) );
  AOI22X1 U71 ( .A0(\d<31> ), .A1(n38), .B0(\q<31> ), .B1(n37), .Y(n79) );
  INVX1 U72 ( .A(n109), .Y(n76) );
  INVX1 U73 ( .A(n108), .Y(n75) );
  INVX1 U74 ( .A(n107), .Y(n74) );
  INVX1 U75 ( .A(n106), .Y(n73) );
  INVX1 U76 ( .A(n105), .Y(n72) );
  INVX1 U77 ( .A(n104), .Y(n71) );
  INVX1 U78 ( .A(n103), .Y(n70) );
  INVXL U79 ( .A(reset), .Y(n78) );
endmodule


module flopr_WIDTH32_0 ( clk, reset, .d({\d<31> , \d<30> , \d<29> , \d<28> , 
        \d<27> , \d<26> , \d<25> , \d<24> , \d<23> , \d<22> , \d<21> , \d<20> , 
        \d<19> , \d<18> , \d<17> , \d<16> , \d<15> , \d<14> , \d<13> , \d<12> , 
        \d<11> , \d<10> , \d<9> , \d<8> , \d<7> , \d<6> , \d<5> , \d<4> , 
        \d<3> , \d<2> , \d<1> , \d<0> }), .q({\q<31> , \q<30> , \q<29> , 
        \q<28> , \q<27> , \q<26> , \q<25> , \q<24> , \q<23> , \q<22> , \q<21> , 
        \q<20> , \q<19> , \q<18> , \q<17> , \q<16> , \q<15> , \q<14> , \q<13> , 
        \q<12> , \q<11> , \q<10> , \q<9> , \q<8> , \q<7> , \q<6> , \q<5> , 
        \q<4> , \q<3> , \q<2> , \q<1> , \q<0> }) );
  input clk, reset, \d<31> , \d<30> , \d<29> , \d<28> , \d<27> , \d<26> ,
         \d<25> , \d<24> , \d<23> , \d<22> , \d<21> , \d<20> , \d<19> ,
         \d<18> , \d<17> , \d<16> , \d<15> , \d<14> , \d<13> , \d<12> ,
         \d<11> , \d<10> , \d<9> , \d<8> , \d<7> , \d<6> , \d<5> , \d<4> ,
         \d<3> , \d<2> , \d<1> , \d<0> ;
  output \q<31> , \q<30> , \q<29> , \q<28> , \q<27> , \q<26> , \q<25> ,
         \q<24> , \q<23> , \q<22> , \q<21> , \q<20> , \q<19> , \q<18> ,
         \q<17> , \q<16> , \q<15> , \q<14> , \q<13> , \q<12> , \q<11> ,
         \q<10> , \q<9> , \q<8> , \q<7> , \q<6> , \q<5> , \q<4> , \q<3> ,
         \q<2> , \q<1> , \q<0> ;
  wire   n1, n2, n3, n4;

  DFFRHQXL \q_reg<31>  ( .D(\d<31> ), .CK(clk), .RN(n1), .Q(\q<31> ) );
  DFFRHQXL \q_reg<30>  ( .D(\d<30> ), .CK(clk), .RN(n1), .Q(\q<30> ) );
  DFFRHQXL \q_reg<29>  ( .D(\d<29> ), .CK(clk), .RN(n1), .Q(\q<29> ) );
  DFFRHQXL \q_reg<28>  ( .D(\d<28> ), .CK(clk), .RN(n1), .Q(\q<28> ) );
  DFFRHQXL \q_reg<27>  ( .D(\d<27> ), .CK(clk), .RN(n1), .Q(\q<27> ) );
  DFFRHQXL \q_reg<26>  ( .D(\d<26> ), .CK(clk), .RN(n1), .Q(\q<26> ) );
  DFFRHQXL \q_reg<25>  ( .D(\d<25> ), .CK(clk), .RN(n1), .Q(\q<25> ) );
  DFFRHQXL \q_reg<24>  ( .D(\d<24> ), .CK(clk), .RN(n1), .Q(\q<24> ) );
  DFFRHQXL \q_reg<23>  ( .D(\d<23> ), .CK(clk), .RN(n1), .Q(\q<23> ) );
  DFFRHQXL \q_reg<22>  ( .D(\d<22> ), .CK(clk), .RN(n1), .Q(\q<22> ) );
  DFFRHQXL \q_reg<21>  ( .D(\d<21> ), .CK(clk), .RN(n1), .Q(\q<21> ) );
  DFFRHQXL \q_reg<20>  ( .D(\d<20> ), .CK(clk), .RN(n1), .Q(\q<20> ) );
  DFFRHQXL \q_reg<19>  ( .D(\d<19> ), .CK(clk), .RN(n2), .Q(\q<19> ) );
  DFFRHQXL \q_reg<18>  ( .D(\d<18> ), .CK(clk), .RN(n2), .Q(\q<18> ) );
  DFFRHQXL \q_reg<17>  ( .D(\d<17> ), .CK(clk), .RN(n2), .Q(\q<17> ) );
  DFFRHQXL \q_reg<16>  ( .D(\d<16> ), .CK(clk), .RN(n2), .Q(\q<16> ) );
  DFFRHQXL \q_reg<15>  ( .D(\d<15> ), .CK(clk), .RN(n2), .Q(\q<15> ) );
  DFFRHQXL \q_reg<14>  ( .D(\d<14> ), .CK(clk), .RN(n2), .Q(\q<14> ) );
  DFFRHQXL \q_reg<13>  ( .D(\d<13> ), .CK(clk), .RN(n2), .Q(\q<13> ) );
  DFFRHQXL \q_reg<12>  ( .D(\d<12> ), .CK(clk), .RN(n2), .Q(\q<12> ) );
  DFFRHQXL \q_reg<11>  ( .D(\d<11> ), .CK(clk), .RN(n2), .Q(\q<11> ) );
  DFFRHQXL \q_reg<10>  ( .D(\d<10> ), .CK(clk), .RN(n2), .Q(\q<10> ) );
  DFFRHQXL \q_reg<9>  ( .D(\d<9> ), .CK(clk), .RN(n2), .Q(\q<9> ) );
  DFFRHQXL \q_reg<8>  ( .D(\d<8> ), .CK(clk), .RN(n2), .Q(\q<8> ) );
  DFFRHQXL \q_reg<7>  ( .D(\d<7> ), .CK(clk), .RN(n1), .Q(\q<7> ) );
  DFFRHQXL \q_reg<6>  ( .D(\d<6> ), .CK(clk), .RN(n2), .Q(\q<6> ) );
  DFFRHQXL \q_reg<5>  ( .D(\d<5> ), .CK(clk), .RN(n1), .Q(\q<5> ) );
  DFFRHQXL \q_reg<4>  ( .D(\d<4> ), .CK(clk), .RN(n2), .Q(\q<4> ) );
  DFFRHQXL \q_reg<3>  ( .D(\d<3> ), .CK(clk), .RN(n1), .Q(\q<3> ) );
  DFFRHQXL \q_reg<2>  ( .D(\d<2> ), .CK(clk), .RN(n2), .Q(\q<2> ) );
  DFFRHQXL \q_reg<1>  ( .D(\d<1> ), .CK(clk), .RN(n4), .Q(\q<1> ) );
  DFFRHQXL \q_reg<0>  ( .D(\d<0> ), .CK(clk), .RN(n4), .Q(\q<0> ) );
  CLKINVX3 U3 ( .A(n3), .Y(n2) );
  CLKINVX3 U4 ( .A(n3), .Y(n1) );
  INVX1 U5 ( .A(n4), .Y(n3) );
  INVXL U6 ( .A(reset), .Y(n4) );
endmodule


module flopr_WIDTH32_3 ( clk, reset, .d({\d<31> , \d<30> , \d<29> , \d<28> , 
        \d<27> , \d<26> , \d<25> , \d<24> , \d<23> , \d<22> , \d<21> , \d<20> , 
        \d<19> , \d<18> , \d<17> , \d<16> , \d<15> , \d<14> , \d<13> , \d<12> , 
        \d<11> , \d<10> , \d<9> , \d<8> , \d<7> , \d<6> , \d<5> , \d<4> , 
        \d<3> , \d<2> , \d<1> , \d<0> }), .q({\q<31> , \q<30> , \q<29> , 
        \q<28> , \q<27> , \q<26> , \q<25> , \q<24> , \q<23> , \q<22> , \q<21> , 
        \q<20> , \q<19> , \q<18> , \q<17> , \q<16> , \q<15> , \q<14> , \q<13> , 
        \q<12> , \q<11> , \q<10> , \q<9> , \q<8> , \q<7> , \q<6> , \q<5> , 
        \q<4> , \q<3> , \q<2> , \q<1> , \q<0> }) );
  input clk, reset, \d<31> , \d<30> , \d<29> , \d<28> , \d<27> , \d<26> ,
         \d<25> , \d<24> , \d<23> , \d<22> , \d<21> , \d<20> , \d<19> ,
         \d<18> , \d<17> , \d<16> , \d<15> , \d<14> , \d<13> , \d<12> ,
         \d<11> , \d<10> , \d<9> , \d<8> , \d<7> , \d<6> , \d<5> , \d<4> ,
         \d<3> , \d<2> , \d<1> , \d<0> ;
  output \q<31> , \q<30> , \q<29> , \q<28> , \q<27> , \q<26> , \q<25> ,
         \q<24> , \q<23> , \q<22> , \q<21> , \q<20> , \q<19> , \q<18> ,
         \q<17> , \q<16> , \q<15> , \q<14> , \q<13> , \q<12> , \q<11> ,
         \q<10> , \q<9> , \q<8> , \q<7> , \q<6> , \q<5> , \q<4> , \q<3> ,
         \q<2> , \q<1> , \q<0> ;
  wire   n1, n2, n3, n4;

  DFFRHQXL \q_reg<31>  ( .D(\d<31> ), .CK(clk), .RN(n1), .Q(\q<31> ) );
  DFFRHQXL \q_reg<30>  ( .D(\d<30> ), .CK(clk), .RN(n1), .Q(\q<30> ) );
  DFFRHQXL \q_reg<29>  ( .D(\d<29> ), .CK(clk), .RN(n1), .Q(\q<29> ) );
  DFFRHQXL \q_reg<28>  ( .D(\d<28> ), .CK(clk), .RN(n1), .Q(\q<28> ) );
  DFFRHQXL \q_reg<27>  ( .D(\d<27> ), .CK(clk), .RN(n1), .Q(\q<27> ) );
  DFFRHQXL \q_reg<26>  ( .D(\d<26> ), .CK(clk), .RN(n1), .Q(\q<26> ) );
  DFFRHQXL \q_reg<25>  ( .D(\d<25> ), .CK(clk), .RN(n1), .Q(\q<25> ) );
  DFFRHQXL \q_reg<24>  ( .D(\d<24> ), .CK(clk), .RN(n1), .Q(\q<24> ) );
  DFFRHQXL \q_reg<23>  ( .D(\d<23> ), .CK(clk), .RN(n1), .Q(\q<23> ) );
  DFFRHQXL \q_reg<22>  ( .D(\d<22> ), .CK(clk), .RN(n1), .Q(\q<22> ) );
  DFFRHQXL \q_reg<21>  ( .D(\d<21> ), .CK(clk), .RN(n1), .Q(\q<21> ) );
  DFFRHQXL \q_reg<20>  ( .D(\d<20> ), .CK(clk), .RN(n1), .Q(\q<20> ) );
  DFFRHQXL \q_reg<19>  ( .D(\d<19> ), .CK(clk), .RN(n2), .Q(\q<19> ) );
  DFFRHQXL \q_reg<18>  ( .D(\d<18> ), .CK(clk), .RN(n2), .Q(\q<18> ) );
  DFFRHQXL \q_reg<17>  ( .D(\d<17> ), .CK(clk), .RN(n2), .Q(\q<17> ) );
  DFFRHQXL \q_reg<16>  ( .D(\d<16> ), .CK(clk), .RN(n2), .Q(\q<16> ) );
  DFFRHQXL \q_reg<15>  ( .D(\d<15> ), .CK(clk), .RN(n2), .Q(\q<15> ) );
  DFFRHQXL \q_reg<14>  ( .D(\d<14> ), .CK(clk), .RN(n2), .Q(\q<14> ) );
  DFFRHQXL \q_reg<13>  ( .D(\d<13> ), .CK(clk), .RN(n2), .Q(\q<13> ) );
  DFFRHQXL \q_reg<12>  ( .D(\d<12> ), .CK(clk), .RN(n2), .Q(\q<12> ) );
  DFFRHQXL \q_reg<11>  ( .D(\d<11> ), .CK(clk), .RN(n2), .Q(\q<11> ) );
  DFFRHQXL \q_reg<10>  ( .D(\d<10> ), .CK(clk), .RN(n2), .Q(\q<10> ) );
  DFFRHQXL \q_reg<9>  ( .D(\d<9> ), .CK(clk), .RN(n2), .Q(\q<9> ) );
  DFFRHQXL \q_reg<8>  ( .D(\d<8> ), .CK(clk), .RN(n2), .Q(\q<8> ) );
  DFFRHQXL \q_reg<7>  ( .D(\d<7> ), .CK(clk), .RN(n1), .Q(\q<7> ) );
  DFFRHQXL \q_reg<6>  ( .D(\d<6> ), .CK(clk), .RN(n2), .Q(\q<6> ) );
  DFFRHQXL \q_reg<5>  ( .D(\d<5> ), .CK(clk), .RN(n1), .Q(\q<5> ) );
  DFFRHQXL \q_reg<4>  ( .D(\d<4> ), .CK(clk), .RN(n2), .Q(\q<4> ) );
  DFFRHQXL \q_reg<3>  ( .D(\d<3> ), .CK(clk), .RN(n1), .Q(\q<3> ) );
  DFFRHQXL \q_reg<2>  ( .D(\d<2> ), .CK(clk), .RN(n2), .Q(\q<2> ) );
  DFFRHQXL \q_reg<1>  ( .D(\d<1> ), .CK(clk), .RN(n4), .Q(\q<1> ) );
  DFFRHQXL \q_reg<0>  ( .D(\d<0> ), .CK(clk), .RN(n4), .Q(\q<0> ) );
  CLKINVX3 U3 ( .A(n3), .Y(n2) );
  CLKINVX3 U4 ( .A(n3), .Y(n1) );
  INVX1 U5 ( .A(n4), .Y(n3) );
  INVXL U6 ( .A(reset), .Y(n4) );
endmodule


module flopr_WIDTH32_2 ( clk, reset, .d({\d<31> , \d<30> , \d<29> , \d<28> , 
        \d<27> , \d<26> , \d<25> , \d<24> , \d<23> , \d<22> , \d<21> , \d<20> , 
        \d<19> , \d<18> , \d<17> , \d<16> , \d<15> , \d<14> , \d<13> , \d<12> , 
        \d<11> , \d<10> , \d<9> , \d<8> , \d<7> , \d<6> , \d<5> , \d<4> , 
        \d<3> , \d<2> , \d<1> , \d<0> }), .q({\q<31> , \q<30> , \q<29> , 
        \q<28> , \q<27> , \q<26> , \q<25> , \q<24> , \q<23> , \q<22> , \q<21> , 
        \q<20> , \q<19> , \q<18> , \q<17> , \q<16> , \q<15> , \q<14> , \q<13> , 
        \q<12> , \q<11> , \q<10> , \q<9> , \q<8> , \q<7> , \q<6> , \q<5> , 
        \q<4> , \q<3> , \q<2> , \q<1> , \q<0> }) );
  input clk, reset, \d<31> , \d<30> , \d<29> , \d<28> , \d<27> , \d<26> ,
         \d<25> , \d<24> , \d<23> , \d<22> , \d<21> , \d<20> , \d<19> ,
         \d<18> , \d<17> , \d<16> , \d<15> , \d<14> , \d<13> , \d<12> ,
         \d<11> , \d<10> , \d<9> , \d<8> , \d<7> , \d<6> , \d<5> , \d<4> ,
         \d<3> , \d<2> , \d<1> , \d<0> ;
  output \q<31> , \q<30> , \q<29> , \q<28> , \q<27> , \q<26> , \q<25> ,
         \q<24> , \q<23> , \q<22> , \q<21> , \q<20> , \q<19> , \q<18> ,
         \q<17> , \q<16> , \q<15> , \q<14> , \q<13> , \q<12> , \q<11> ,
         \q<10> , \q<9> , \q<8> , \q<7> , \q<6> , \q<5> , \q<4> , \q<3> ,
         \q<2> , \q<1> , \q<0> ;
  wire   n1, n2, n3, n4;

  DFFRHQXL \q_reg<31>  ( .D(\d<31> ), .CK(clk), .RN(n1), .Q(\q<31> ) );
  DFFRHQXL \q_reg<30>  ( .D(\d<30> ), .CK(clk), .RN(n1), .Q(\q<30> ) );
  DFFRHQXL \q_reg<29>  ( .D(\d<29> ), .CK(clk), .RN(n1), .Q(\q<29> ) );
  DFFRHQXL \q_reg<28>  ( .D(\d<28> ), .CK(clk), .RN(n1), .Q(\q<28> ) );
  DFFRHQXL \q_reg<27>  ( .D(\d<27> ), .CK(clk), .RN(n1), .Q(\q<27> ) );
  DFFRHQXL \q_reg<26>  ( .D(\d<26> ), .CK(clk), .RN(n1), .Q(\q<26> ) );
  DFFRHQXL \q_reg<25>  ( .D(\d<25> ), .CK(clk), .RN(n1), .Q(\q<25> ) );
  DFFRHQXL \q_reg<24>  ( .D(\d<24> ), .CK(clk), .RN(n1), .Q(\q<24> ) );
  DFFRHQXL \q_reg<23>  ( .D(\d<23> ), .CK(clk), .RN(n1), .Q(\q<23> ) );
  DFFRHQXL \q_reg<22>  ( .D(\d<22> ), .CK(clk), .RN(n1), .Q(\q<22> ) );
  DFFRHQXL \q_reg<21>  ( .D(\d<21> ), .CK(clk), .RN(n1), .Q(\q<21> ) );
  DFFRHQXL \q_reg<20>  ( .D(\d<20> ), .CK(clk), .RN(n1), .Q(\q<20> ) );
  DFFRHQXL \q_reg<19>  ( .D(\d<19> ), .CK(clk), .RN(n2), .Q(\q<19> ) );
  DFFRHQXL \q_reg<18>  ( .D(\d<18> ), .CK(clk), .RN(n2), .Q(\q<18> ) );
  DFFRHQXL \q_reg<17>  ( .D(\d<17> ), .CK(clk), .RN(n2), .Q(\q<17> ) );
  DFFRHQXL \q_reg<16>  ( .D(\d<16> ), .CK(clk), .RN(n2), .Q(\q<16> ) );
  DFFRHQXL \q_reg<15>  ( .D(\d<15> ), .CK(clk), .RN(n2), .Q(\q<15> ) );
  DFFRHQXL \q_reg<14>  ( .D(\d<14> ), .CK(clk), .RN(n2), .Q(\q<14> ) );
  DFFRHQXL \q_reg<13>  ( .D(\d<13> ), .CK(clk), .RN(n2), .Q(\q<13> ) );
  DFFRHQXL \q_reg<12>  ( .D(\d<12> ), .CK(clk), .RN(n2), .Q(\q<12> ) );
  DFFRHQXL \q_reg<11>  ( .D(\d<11> ), .CK(clk), .RN(n2), .Q(\q<11> ) );
  DFFRHQXL \q_reg<10>  ( .D(\d<10> ), .CK(clk), .RN(n2), .Q(\q<10> ) );
  DFFRHQXL \q_reg<9>  ( .D(\d<9> ), .CK(clk), .RN(n2), .Q(\q<9> ) );
  DFFRHQXL \q_reg<8>  ( .D(\d<8> ), .CK(clk), .RN(n2), .Q(\q<8> ) );
  DFFRHQXL \q_reg<7>  ( .D(\d<7> ), .CK(clk), .RN(n1), .Q(\q<7> ) );
  DFFRHQXL \q_reg<6>  ( .D(\d<6> ), .CK(clk), .RN(n2), .Q(\q<6> ) );
  DFFRHQXL \q_reg<5>  ( .D(\d<5> ), .CK(clk), .RN(n1), .Q(\q<5> ) );
  DFFRHQXL \q_reg<4>  ( .D(\d<4> ), .CK(clk), .RN(n2), .Q(\q<4> ) );
  DFFRHQXL \q_reg<3>  ( .D(\d<3> ), .CK(clk), .RN(n1), .Q(\q<3> ) );
  DFFRHQXL \q_reg<2>  ( .D(\d<2> ), .CK(clk), .RN(n2), .Q(\q<2> ) );
  DFFRHQXL \q_reg<1>  ( .D(\d<1> ), .CK(clk), .RN(n4), .Q(\q<1> ) );
  DFFRHQXL \q_reg<0>  ( .D(\d<0> ), .CK(clk), .RN(n4), .Q(\q<0> ) );
  CLKINVX3 U3 ( .A(n3), .Y(n2) );
  CLKINVX3 U4 ( .A(n3), .Y(n1) );
  INVX1 U5 ( .A(n4), .Y(n3) );
  INVXL U6 ( .A(reset), .Y(n4) );
endmodule


module flopr_WIDTH32_1 ( clk, reset, .d({\d<31> , \d<30> , \d<29> , \d<28> , 
        \d<27> , \d<26> , \d<25> , \d<24> , \d<23> , \d<22> , \d<21> , \d<20> , 
        \d<19> , \d<18> , \d<17> , \d<16> , \d<15> , \d<14> , \d<13> , \d<12> , 
        \d<11> , \d<10> , \d<9> , \d<8> , \d<7> , \d<6> , \d<5> , \d<4> , 
        \d<3> , \d<2> , \d<1> , \d<0> }), .q({\q<31> , \q<30> , \q<29> , 
        \q<28> , \q<27> , \q<26> , \q<25> , \q<24> , \q<23> , \q<22> , \q<21> , 
        \q<20> , \q<19> , \q<18> , \q<17> , \q<16> , \q<15> , \q<14> , \q<13> , 
        \q<12> , \q<11> , \q<10> , \q<9> , \q<8> , \q<7> , \q<6> , \q<5> , 
        \q<4> , \q<3> , \q<2> , \q<1> , \q<0> }) );
  input clk, reset, \d<31> , \d<30> , \d<29> , \d<28> , \d<27> , \d<26> ,
         \d<25> , \d<24> , \d<23> , \d<22> , \d<21> , \d<20> , \d<19> ,
         \d<18> , \d<17> , \d<16> , \d<15> , \d<14> , \d<13> , \d<12> ,
         \d<11> , \d<10> , \d<9> , \d<8> , \d<7> , \d<6> , \d<5> , \d<4> ,
         \d<3> , \d<2> , \d<1> , \d<0> ;
  output \q<31> , \q<30> , \q<29> , \q<28> , \q<27> , \q<26> , \q<25> ,
         \q<24> , \q<23> , \q<22> , \q<21> , \q<20> , \q<19> , \q<18> ,
         \q<17> , \q<16> , \q<15> , \q<14> , \q<13> , \q<12> , \q<11> ,
         \q<10> , \q<9> , \q<8> , \q<7> , \q<6> , \q<5> , \q<4> , \q<3> ,
         \q<2> , \q<1> , \q<0> ;
  wire   n1, n2, n3, n4;

  DFFRHQXL \q_reg<31>  ( .D(\d<31> ), .CK(clk), .RN(n1), .Q(\q<31> ) );
  DFFRHQXL \q_reg<30>  ( .D(\d<30> ), .CK(clk), .RN(n1), .Q(\q<30> ) );
  DFFRHQXL \q_reg<29>  ( .D(\d<29> ), .CK(clk), .RN(n1), .Q(\q<29> ) );
  DFFRHQXL \q_reg<28>  ( .D(\d<28> ), .CK(clk), .RN(n1), .Q(\q<28> ) );
  DFFRHQXL \q_reg<27>  ( .D(\d<27> ), .CK(clk), .RN(n1), .Q(\q<27> ) );
  DFFRHQXL \q_reg<26>  ( .D(\d<26> ), .CK(clk), .RN(n1), .Q(\q<26> ) );
  DFFRHQXL \q_reg<25>  ( .D(\d<25> ), .CK(clk), .RN(n1), .Q(\q<25> ) );
  DFFRHQXL \q_reg<24>  ( .D(\d<24> ), .CK(clk), .RN(n1), .Q(\q<24> ) );
  DFFRHQXL \q_reg<23>  ( .D(\d<23> ), .CK(clk), .RN(n1), .Q(\q<23> ) );
  DFFRHQXL \q_reg<22>  ( .D(\d<22> ), .CK(clk), .RN(n1), .Q(\q<22> ) );
  DFFRHQXL \q_reg<21>  ( .D(\d<21> ), .CK(clk), .RN(n1), .Q(\q<21> ) );
  DFFRHQXL \q_reg<20>  ( .D(\d<20> ), .CK(clk), .RN(n1), .Q(\q<20> ) );
  DFFRHQXL \q_reg<19>  ( .D(\d<19> ), .CK(clk), .RN(n2), .Q(\q<19> ) );
  DFFRHQXL \q_reg<18>  ( .D(\d<18> ), .CK(clk), .RN(n2), .Q(\q<18> ) );
  DFFRHQXL \q_reg<17>  ( .D(\d<17> ), .CK(clk), .RN(n2), .Q(\q<17> ) );
  DFFRHQXL \q_reg<16>  ( .D(\d<16> ), .CK(clk), .RN(n2), .Q(\q<16> ) );
  DFFRHQXL \q_reg<15>  ( .D(\d<15> ), .CK(clk), .RN(n2), .Q(\q<15> ) );
  DFFRHQXL \q_reg<14>  ( .D(\d<14> ), .CK(clk), .RN(n2), .Q(\q<14> ) );
  DFFRHQXL \q_reg<13>  ( .D(\d<13> ), .CK(clk), .RN(n2), .Q(\q<13> ) );
  DFFRHQXL \q_reg<12>  ( .D(\d<12> ), .CK(clk), .RN(n2), .Q(\q<12> ) );
  DFFRHQXL \q_reg<9>  ( .D(\d<9> ), .CK(clk), .RN(n2), .Q(\q<9> ) );
  DFFRHQXL \q_reg<11>  ( .D(\d<11> ), .CK(clk), .RN(n2), .Q(\q<11> ) );
  DFFRHQXL \q_reg<10>  ( .D(\d<10> ), .CK(clk), .RN(n2), .Q(\q<10> ) );
  DFFRHQXL \q_reg<8>  ( .D(\d<8> ), .CK(clk), .RN(n2), .Q(\q<8> ) );
  DFFRHQXL \q_reg<7>  ( .D(\d<7> ), .CK(clk), .RN(n1), .Q(\q<7> ) );
  DFFRHQXL \q_reg<6>  ( .D(\d<6> ), .CK(clk), .RN(n2), .Q(\q<6> ) );
  DFFRHQXL \q_reg<5>  ( .D(\d<5> ), .CK(clk), .RN(n1), .Q(\q<5> ) );
  DFFRHQXL \q_reg<4>  ( .D(\d<4> ), .CK(clk), .RN(n2), .Q(\q<4> ) );
  DFFRHQXL \q_reg<3>  ( .D(\d<3> ), .CK(clk), .RN(n1), .Q(\q<3> ) );
  DFFRHQXL \q_reg<2>  ( .D(\d<2> ), .CK(clk), .RN(n2), .Q(\q<2> ) );
  DFFRHQXL \q_reg<1>  ( .D(\d<1> ), .CK(clk), .RN(n4), .Q(\q<1> ) );
  DFFRHQXL \q_reg<0>  ( .D(\d<0> ), .CK(clk), .RN(n4), .Q(\q<0> ) );
  CLKINVX3 U3 ( .A(n3), .Y(n2) );
  CLKINVX3 U4 ( .A(n3), .Y(n1) );
  INVX1 U5 ( .A(n4), .Y(n3) );
  INVXL U6 ( .A(reset), .Y(n4) );
endmodule


module mux2_WIDTH32 ( .d0({\d0<31> , \d0<30> , \d0<29> , \d0<28> , \d0<27> , 
        \d0<26> , \d0<25> , \d0<24> , \d0<23> , \d0<22> , \d0<21> , \d0<20> , 
        \d0<19> , \d0<18> , \d0<17> , \d0<16> , \d0<15> , \d0<14> , \d0<13> , 
        \d0<12> , \d0<11> , \d0<10> , \d0<9> , \d0<8> , \d0<7> , \d0<6> , 
        \d0<5> , \d0<4> , \d0<3> , \d0<2> , \d0<1> , \d0<0> }), .d1({\d1<31> , 
        \d1<30> , \d1<29> , \d1<28> , \d1<27> , \d1<26> , \d1<25> , \d1<24> , 
        \d1<23> , \d1<22> , \d1<21> , \d1<20> , \d1<19> , \d1<18> , \d1<17> , 
        \d1<16> , \d1<15> , \d1<14> , \d1<13> , \d1<12> , \d1<11> , \d1<10> , 
        \d1<9> , \d1<8> , \d1<7> , \d1<6> , \d1<5> , \d1<4> , \d1<3> , \d1<2> , 
        \d1<1> , \d1<0> }), s, .y({\y<31> , \y<30> , \y<29> , \y<28> , \y<27> , 
        \y<26> , \y<25> , \y<24> , \y<23> , \y<22> , \y<21> , \y<20> , \y<19> , 
        \y<18> , \y<17> , \y<16> , \y<15> , \y<14> , \y<13> , \y<12> , \y<11> , 
        \y<10> , \y<9> , \y<8> , \y<7> , \y<6> , \y<5> , \y<4> , \y<3> , 
        \y<2> , \y<1> , \y<0> }) );
  input \d0<31> , \d0<30> , \d0<29> , \d0<28> , \d0<27> , \d0<26> , \d0<25> ,
         \d0<24> , \d0<23> , \d0<22> , \d0<21> , \d0<20> , \d0<19> , \d0<18> ,
         \d0<17> , \d0<16> , \d0<15> , \d0<14> , \d0<13> , \d0<12> , \d0<11> ,
         \d0<10> , \d0<9> , \d0<8> , \d0<7> , \d0<6> , \d0<5> , \d0<4> ,
         \d0<3> , \d0<2> , \d0<1> , \d0<0> , \d1<31> , \d1<30> , \d1<29> ,
         \d1<28> , \d1<27> , \d1<26> , \d1<25> , \d1<24> , \d1<23> , \d1<22> ,
         \d1<21> , \d1<20> , \d1<19> , \d1<18> , \d1<17> , \d1<16> , \d1<15> ,
         \d1<14> , \d1<13> , \d1<12> , \d1<11> , \d1<10> , \d1<9> , \d1<8> ,
         \d1<7> , \d1<6> , \d1<5> , \d1<4> , \d1<3> , \d1<2> , \d1<1> ,
         \d1<0> , s;
  output \y<31> , \y<30> , \y<29> , \y<28> , \y<27> , \y<26> , \y<25> ,
         \y<24> , \y<23> , \y<22> , \y<21> , \y<20> , \y<19> , \y<18> ,
         \y<17> , \y<16> , \y<15> , \y<14> , \y<13> , \y<12> , \y<11> ,
         \y<10> , \y<9> , \y<8> , \y<7> , \y<6> , \y<5> , \y<4> , \y<3> ,
         \y<2> , \y<1> , \y<0> ;
  wire   n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62,
         n63, n64, n65, n66, n1, n2, n3, n4, n5, n6, n7;

  AOI22XL U1 ( .A0(\d0<0> ), .A1(n1), .B0(\d1<0> ), .B1(n6), .Y(n66) );
  AOI22XL U2 ( .A0(\d0<1> ), .A1(n1), .B0(\d1<1> ), .B1(n3), .Y(n55) );
  AOI22XL U3 ( .A0(\d0<2> ), .A1(n2), .B0(\d1<2> ), .B1(n4), .Y(n44) );
  AOI22XL U4 ( .A0(\d0<3> ), .A1(n2), .B0(\d1<3> ), .B1(n4), .Y(n41) );
  AOI22XL U5 ( .A0(\d0<4> ), .A1(n1), .B0(\d1<4> ), .B1(n6), .Y(n40) );
  AOI22XL U6 ( .A0(\d0<5> ), .A1(n2), .B0(\d1<5> ), .B1(n3), .Y(n39) );
  AOI22XL U7 ( .A0(\d0<6> ), .A1(n1), .B0(\d1<6> ), .B1(n3), .Y(n38) );
  AOI22XL U8 ( .A0(\d0<7> ), .A1(n2), .B0(\d1<7> ), .B1(n4), .Y(n37) );
  AOI22XL U9 ( .A0(\d0<8> ), .A1(n1), .B0(\d1<8> ), .B1(n3), .Y(n36) );
  AOI22XL U10 ( .A0(\d0<9> ), .A1(n7), .B0(n6), .B1(\d1<9> ), .Y(n35) );
  AOI22XL U11 ( .A0(\d0<10> ), .A1(n1), .B0(\d1<10> ), .B1(n5), .Y(n65) );
  AOI22XL U12 ( .A0(\d0<11> ), .A1(n1), .B0(\d1<11> ), .B1(s), .Y(n64) );
  AOI22XL U13 ( .A0(\d0<12> ), .A1(n1), .B0(\d1<12> ), .B1(n4), .Y(n63) );
  AOI22XL U14 ( .A0(\d0<13> ), .A1(n1), .B0(\d1<13> ), .B1(n6), .Y(n62) );
  AOI22XL U15 ( .A0(\d0<14> ), .A1(n1), .B0(\d1<14> ), .B1(n3), .Y(n61) );
  AOI22XL U16 ( .A0(\d0<15> ), .A1(n1), .B0(\d1<15> ), .B1(n6), .Y(n60) );
  AOI22XL U17 ( .A0(\d0<16> ), .A1(n1), .B0(\d1<16> ), .B1(s), .Y(n59) );
  AOI22XL U18 ( .A0(\d0<17> ), .A1(n1), .B0(\d1<17> ), .B1(n6), .Y(n58) );
  AOI22XL U19 ( .A0(\d0<18> ), .A1(n1), .B0(\d1<18> ), .B1(n4), .Y(n57) );
  AOI22XL U20 ( .A0(\d0<19> ), .A1(n1), .B0(\d1<19> ), .B1(n3), .Y(n56) );
  AOI22XL U21 ( .A0(\d0<20> ), .A1(n2), .B0(\d1<20> ), .B1(n5), .Y(n54) );
  AOI22XL U22 ( .A0(\d0<21> ), .A1(n2), .B0(\d1<21> ), .B1(s), .Y(n53) );
  AOI22XL U23 ( .A0(\d0<22> ), .A1(n2), .B0(\d1<22> ), .B1(n5), .Y(n52) );
  AOI22XL U24 ( .A0(\d0<23> ), .A1(n2), .B0(\d1<23> ), .B1(n5), .Y(n51) );
  AOI22XL U25 ( .A0(\d0<24> ), .A1(n2), .B0(\d1<24> ), .B1(n6), .Y(n50) );
  AOI22XL U26 ( .A0(\d0<25> ), .A1(n2), .B0(\d1<25> ), .B1(s), .Y(n49) );
  AOI22XL U27 ( .A0(\d0<26> ), .A1(n2), .B0(\d1<26> ), .B1(s), .Y(n48) );
  AOI22XL U28 ( .A0(\d0<27> ), .A1(n2), .B0(\d1<27> ), .B1(s), .Y(n47) );
  AOI22XL U29 ( .A0(\d0<28> ), .A1(n2), .B0(\d1<28> ), .B1(n5), .Y(n46) );
  AOI22XL U30 ( .A0(\d0<29> ), .A1(n2), .B0(\d1<29> ), .B1(n4), .Y(n45) );
  AOI22XL U31 ( .A0(\d0<30> ), .A1(n2), .B0(\d1<30> ), .B1(n5), .Y(n43) );
  CLKINVX3 U32 ( .A(n5), .Y(n1) );
  CLKINVX3 U33 ( .A(n3), .Y(n2) );
  INVX1 U34 ( .A(n7), .Y(n3) );
  INVX1 U35 ( .A(n7), .Y(n5) );
  INVX1 U36 ( .A(n7), .Y(n4) );
  INVX1 U37 ( .A(n7), .Y(n6) );
  INVX1 U38 ( .A(s), .Y(n7) );
  INVX1 U39 ( .A(n35), .Y(\y<9> ) );
  INVX1 U40 ( .A(n66), .Y(\y<0> ) );
  INVX1 U41 ( .A(n55), .Y(\y<1> ) );
  INVX1 U42 ( .A(n44), .Y(\y<2> ) );
  INVX1 U43 ( .A(n65), .Y(\y<10> ) );
  INVX1 U44 ( .A(n64), .Y(\y<11> ) );
  INVX1 U45 ( .A(n63), .Y(\y<12> ) );
  INVX1 U46 ( .A(n62), .Y(\y<13> ) );
  INVX1 U47 ( .A(n61), .Y(\y<14> ) );
  INVX1 U48 ( .A(n60), .Y(\y<15> ) );
  INVX1 U49 ( .A(n59), .Y(\y<16> ) );
  INVX1 U50 ( .A(n58), .Y(\y<17> ) );
  INVX1 U51 ( .A(n57), .Y(\y<18> ) );
  INVX1 U52 ( .A(n56), .Y(\y<19> ) );
  INVX1 U53 ( .A(n54), .Y(\y<20> ) );
  INVX1 U54 ( .A(n53), .Y(\y<21> ) );
  INVX1 U55 ( .A(n52), .Y(\y<22> ) );
  INVX1 U56 ( .A(n51), .Y(\y<23> ) );
  INVX1 U57 ( .A(n50), .Y(\y<24> ) );
  INVX1 U58 ( .A(n49), .Y(\y<25> ) );
  INVX1 U59 ( .A(n48), .Y(\y<26> ) );
  INVX1 U60 ( .A(n47), .Y(\y<27> ) );
  INVX1 U61 ( .A(n46), .Y(\y<28> ) );
  INVX1 U62 ( .A(n45), .Y(\y<29> ) );
  INVX1 U63 ( .A(n43), .Y(\y<30> ) );
  INVX1 U64 ( .A(n41), .Y(\y<3> ) );
  INVX1 U65 ( .A(n40), .Y(\y<4> ) );
  INVX1 U66 ( .A(n39), .Y(\y<5> ) );
  INVX1 U67 ( .A(n38), .Y(\y<6> ) );
  INVX1 U68 ( .A(n37), .Y(\y<7> ) );
  INVX1 U69 ( .A(n36), .Y(\y<8> ) );
  INVX1 U70 ( .A(n42), .Y(\y<31> ) );
  AOI22X1 U71 ( .A0(\d0<31> ), .A1(n7), .B0(\d1<31> ), .B1(n4), .Y(n42) );
endmodule


module mux2_WIDTH4_0 ( .d0({\d0<3> , \d0<2> , \d0<1> , \d0<0> }), .d1({\d1<3> , 
        \d1<2> , \d1<1> , \d1<0> }), s, .y({\y<3> , \y<2> , \y<1> , \y<0> })
 );
  input \d0<3> , \d0<2> , \d0<1> , \d0<0> , \d1<3> , \d1<2> , \d1<1> , \d1<0> ,
         s;
  output \y<3> , \y<2> , \y<1> , \y<0> ;
  wire   n7, n8, n9, n10, n1;

  INVX1 U1 ( .A(s), .Y(n1) );
  INVX1 U2 ( .A(n10), .Y(\y<0> ) );
  AOI22X1 U3 ( .A0(\d0<0> ), .A1(n1), .B0(\d1<0> ), .B1(s), .Y(n10) );
  INVX1 U4 ( .A(n7), .Y(\y<3> ) );
  AOI22X1 U5 ( .A0(\d0<3> ), .A1(n1), .B0(s), .B1(\d1<3> ), .Y(n7) );
  INVX1 U6 ( .A(n9), .Y(\y<1> ) );
  AOI22X1 U7 ( .A0(\d0<1> ), .A1(n1), .B0(\d1<1> ), .B1(s), .Y(n9) );
  INVX1 U8 ( .A(n8), .Y(\y<2> ) );
  AOI22X1 U9 ( .A0(\d0<2> ), .A1(n1), .B0(\d1<2> ), .B1(s), .Y(n8) );
endmodule


module mux2_WIDTH4_1 ( .d0({\d0<3> , \d0<2> , \d0<1> , \d0<0> }), .d1({\d1<3> , 
        \d1<2> , \d1<1> , \d1<0> }), s, .y({\y<3> , \y<2> , \y<1> , \y<0> })
 );
  input \d0<3> , \d0<2> , \d0<1> , \d0<0> , \d1<3> , \d1<2> , \d1<1> , \d1<0> ,
         s;
  output \y<3> , \y<2> , \y<1> , \y<0> ;
  wire   n1, n2, n3, n4, n5;

  AOI22XL U1 ( .A0(\d0<0> ), .A1(n1), .B0(\d1<0> ), .B1(s), .Y(n2) );
  AOI22XL U2 ( .A0(\d0<1> ), .A1(n1), .B0(\d1<1> ), .B1(s), .Y(n3) );
  AOI22XL U3 ( .A0(\d0<3> ), .A1(n1), .B0(s), .B1(\d1<3> ), .Y(n5) );
  AOI22XL U4 ( .A0(\d0<2> ), .A1(n1), .B0(\d1<2> ), .B1(s), .Y(n4) );
  INVX1 U5 ( .A(s), .Y(n1) );
  INVX1 U6 ( .A(n2), .Y(\y<0> ) );
  INVX1 U7 ( .A(n3), .Y(\y<1> ) );
  INVX1 U8 ( .A(n4), .Y(\y<2> ) );
  INVX1 U9 ( .A(n5), .Y(\y<3> ) );
endmodule


module mux3_WIDTH32_0 ( .d0({\d0<31> , \d0<30> , \d0<29> , \d0<28> , \d0<27> , 
        \d0<26> , \d0<25> , \d0<24> , \d0<23> , \d0<22> , \d0<21> , \d0<20> , 
        \d0<19> , \d0<18> , \d0<17> , \d0<16> , \d0<15> , \d0<14> , \d0<13> , 
        \d0<12> , \d0<11> , \d0<10> , \d0<9> , \d0<8> , \d0<7> , \d0<6> , 
        \d0<5> , \d0<4> , \d0<3> , \d0<2> , \d0<1> , \d0<0> }), .d1({\d1<31> , 
        \d1<30> , \d1<29> , \d1<28> , \d1<27> , \d1<26> , \d1<25> , \d1<24> , 
        \d1<23> , \d1<22> , \d1<21> , \d1<20> , \d1<19> , \d1<18> , \d1<17> , 
        \d1<16> , \d1<15> , \d1<14> , \d1<13> , \d1<12> , \d1<11> , \d1<10> , 
        \d1<9> , \d1<8> , \d1<7> , \d1<6> , \d1<5> , \d1<4> , \d1<3> , \d1<2> , 
        \d1<1> , \d1<0> }), .d2({\d2<31> , \d2<30> , \d2<29> , \d2<28> , 
        \d2<27> , \d2<26> , \d2<25> , \d2<24> , \d2<23> , \d2<22> , \d2<21> , 
        \d2<20> , \d2<19> , \d2<18> , \d2<17> , \d2<16> , \d2<15> , \d2<14> , 
        \d2<13> , \d2<12> , \d2<11> , \d2<10> , \d2<9> , \d2<8> , \d2<7> , 
        \d2<6> , \d2<5> , \d2<4> , \d2<3> , \d2<2> , \d2<1> , \d2<0> }), .s({
        \s<1> , \s<0> }), .y({\y<31> , \y<30> , \y<29> , \y<28> , \y<27> , 
        \y<26> , \y<25> , \y<24> , \y<23> , \y<22> , \y<21> , \y<20> , \y<19> , 
        \y<18> , \y<17> , \y<16> , \y<15> , \y<14> , \y<13> , \y<12> , \y<11> , 
        \y<10> , \y<9> , \y<8> , \y<7> , \y<6> , \y<5> , \y<4> , \y<3> , 
        \y<2> , \y<1> , \y<0> }) );
  input \d0<31> , \d0<30> , \d0<29> , \d0<28> , \d0<27> , \d0<26> , \d0<25> ,
         \d0<24> , \d0<23> , \d0<22> , \d0<21> , \d0<20> , \d0<19> , \d0<18> ,
         \d0<17> , \d0<16> , \d0<15> , \d0<14> , \d0<13> , \d0<12> , \d0<11> ,
         \d0<10> , \d0<9> , \d0<8> , \d0<7> , \d0<6> , \d0<5> , \d0<4> ,
         \d0<3> , \d0<2> , \d0<1> , \d0<0> , \d1<31> , \d1<30> , \d1<29> ,
         \d1<28> , \d1<27> , \d1<26> , \d1<25> , \d1<24> , \d1<23> , \d1<22> ,
         \d1<21> , \d1<20> , \d1<19> , \d1<18> , \d1<17> , \d1<16> , \d1<15> ,
         \d1<14> , \d1<13> , \d1<12> , \d1<11> , \d1<10> , \d1<9> , \d1<8> ,
         \d1<7> , \d1<6> , \d1<5> , \d1<4> , \d1<3> , \d1<2> , \d1<1> ,
         \d1<0> , \d2<31> , \d2<30> , \d2<29> , \d2<28> , \d2<27> , \d2<26> ,
         \d2<25> , \d2<24> , \d2<23> , \d2<22> , \d2<21> , \d2<20> , \d2<19> ,
         \d2<18> , \d2<17> , \d2<16> , \d2<15> , \d2<14> , \d2<13> , \d2<12> ,
         \d2<11> , \d2<10> , \d2<9> , \d2<8> , \d2<7> , \d2<6> , \d2<5> ,
         \d2<4> , \d2<3> , \d2<2> , \d2<1> , \d2<0> , \s<1> , \s<0> ;
  output \y<31> , \y<30> , \y<29> , \y<28> , \y<27> , \y<26> , \y<25> ,
         \y<24> , \y<23> , \y<22> , \y<21> , \y<20> , \y<19> , \y<18> ,
         \y<17> , \y<16> , \y<15> , \y<14> , \y<13> , \y<12> , \y<11> ,
         \y<10> , \y<9> , \y<8> , \y<7> , \y<6> , \y<5> , \y<4> , \y<3> ,
         \y<2> , \y<1> , \y<0> ;
  wire   n2, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n1, n3, n36, n37, n38, n39, n40, n41, n42;

  BUFX20 U1 ( .A(n38), .Y(n1) );
  BUFX20 U2 ( .A(n4), .Y(n3) );
  BUFX20 U3 ( .A(n1), .Y(n36) );
  OAI2BB1X2 U4 ( .A0N(\d2<0> ), .A1N(n41), .B0(n35), .Y(\y<0> ) );
  BUFX20 U5 ( .A(n1), .Y(n37) );
  NOR2X4 U6 ( .A(\s<0> ), .B(n41), .Y(n38) );
  CLKINVX20 U7 ( .A(n42), .Y(n41) );
  INVX8 U8 ( .A(n40), .Y(n39) );
  OAI2BB1X2 U9 ( .A0N(\d2<2> ), .A1N(n41), .B0(n13), .Y(\y<2> ) );
  OAI2BB1X1 U10 ( .A0N(\d2<3> ), .A1N(n41), .B0(n10), .Y(\y<3> ) );
  OAI2BB1X1 U11 ( .A0N(\d2<4> ), .A1N(n41), .B0(n9), .Y(\y<4> ) );
  AOI22X2 U12 ( .A0(\d0<1> ), .A1(n1), .B0(\d1<1> ), .B1(n3), .Y(n24) );
  AOI22X4 U13 ( .A0(\d0<0> ), .A1(n1), .B0(\d1<0> ), .B1(n3), .Y(n35) );
  AOI22XL U14 ( .A0(\d0<10> ), .A1(n37), .B0(\d1<10> ), .B1(n39), .Y(n34) );
  AOI22XL U15 ( .A0(\d0<11> ), .A1(n36), .B0(\d1<11> ), .B1(n39), .Y(n33) );
  AOI22XL U16 ( .A0(\d0<12> ), .A1(n37), .B0(\d1<12> ), .B1(n39), .Y(n32) );
  OAI2BB1X4 U17 ( .A0N(\d2<1> ), .A1N(n41), .B0(n24), .Y(\y<1> ) );
  AOI22X2 U18 ( .A0(\d0<2> ), .A1(n36), .B0(\d1<2> ), .B1(n3), .Y(n13) );
  NOR2BX4 U19 ( .AN(\s<0> ), .B(n41), .Y(n4) );
  AOI22XL U20 ( .A0(\d0<15> ), .A1(n36), .B0(\d1<15> ), .B1(n39), .Y(n29) );
  AOI22XL U21 ( .A0(\d0<14> ), .A1(n37), .B0(\d1<14> ), .B1(n39), .Y(n30) );
  AOI22XL U22 ( .A0(\d0<13> ), .A1(n36), .B0(\d1<13> ), .B1(n39), .Y(n31) );
  AOI22XL U23 ( .A0(\d0<18> ), .A1(n36), .B0(\d1<18> ), .B1(n39), .Y(n26) );
  AOI22XL U24 ( .A0(\d0<17> ), .A1(n37), .B0(\d1<17> ), .B1(n39), .Y(n27) );
  AOI22XL U25 ( .A0(\d0<16> ), .A1(n37), .B0(\d1<16> ), .B1(n39), .Y(n28) );
  AOI22XL U26 ( .A0(\d0<22> ), .A1(n36), .B0(\d1<22> ), .B1(n39), .Y(n21) );
  AOI22XL U27 ( .A0(\d0<21> ), .A1(n37), .B0(\d1<21> ), .B1(n39), .Y(n22) );
  AOI22XL U28 ( .A0(\d0<20> ), .A1(n36), .B0(\d1<20> ), .B1(n39), .Y(n23) );
  AOI22XL U29 ( .A0(\d0<19> ), .A1(n37), .B0(\d1<19> ), .B1(n39), .Y(n25) );
  AOI22XL U30 ( .A0(\d0<24> ), .A1(n37), .B0(\d1<24> ), .B1(n39), .Y(n19) );
  AOI22XL U31 ( .A0(\d0<23> ), .A1(n37), .B0(\d1<23> ), .B1(n39), .Y(n20) );
  AOI22XL U32 ( .A0(\d0<25> ), .A1(n36), .B0(\d1<25> ), .B1(n39), .Y(n18) );
  AOI22XL U33 ( .A0(\d0<26> ), .A1(n37), .B0(\d1<26> ), .B1(n39), .Y(n17) );
  AOI22XL U34 ( .A0(\d0<27> ), .A1(n36), .B0(\d1<27> ), .B1(n39), .Y(n16) );
  AOI22XL U35 ( .A0(\d0<28> ), .A1(n36), .B0(\d1<28> ), .B1(n39), .Y(n15) );
  AOI22XL U36 ( .A0(\d0<29> ), .A1(n36), .B0(\d1<29> ), .B1(n3), .Y(n14) );
  AOI22XL U37 ( .A0(\d0<30> ), .A1(n37), .B0(\d1<30> ), .B1(n3), .Y(n12) );
  OAI2BB1X1 U38 ( .A0N(\d2<31> ), .A1N(n41), .B0(n11), .Y(\y<31> ) );
  AOI22XL U39 ( .A0(\d0<31> ), .A1(n37), .B0(\d1<31> ), .B1(n39), .Y(n11) );
  INVX1 U40 ( .A(n3), .Y(n40) );
  INVX1 U41 ( .A(\s<1> ), .Y(n42) );
  AOI22X1 U42 ( .A0(\d0<3> ), .A1(n37), .B0(\d1<3> ), .B1(n3), .Y(n10) );
  AOI22X1 U43 ( .A0(\d0<4> ), .A1(n37), .B0(\d1<4> ), .B1(n3), .Y(n9) );
  OAI2BB1X1 U44 ( .A0N(\d2<5> ), .A1N(n41), .B0(n8), .Y(\y<5> ) );
  AOI22X1 U45 ( .A0(\d0<5> ), .A1(n37), .B0(\d1<5> ), .B1(n3), .Y(n8) );
  OAI2BB1X1 U46 ( .A0N(n41), .A1N(\d2<9> ), .B0(n2), .Y(\y<9> ) );
  AOI22X1 U47 ( .A0(\d0<9> ), .A1(n36), .B0(\d1<9> ), .B1(n39), .Y(n2) );
  OAI2BB1X1 U48 ( .A0N(\d2<6> ), .A1N(n41), .B0(n7), .Y(\y<6> ) );
  AOI22X1 U49 ( .A0(\d0<6> ), .A1(n37), .B0(\d1<6> ), .B1(n39), .Y(n7) );
  OAI2BB1X1 U50 ( .A0N(\d2<7> ), .A1N(n41), .B0(n6), .Y(\y<7> ) );
  AOI22X1 U51 ( .A0(\d0<7> ), .A1(n37), .B0(\d1<7> ), .B1(n39), .Y(n6) );
  OAI2BB1X1 U52 ( .A0N(\d2<8> ), .A1N(n41), .B0(n5), .Y(\y<8> ) );
  AOI22X1 U53 ( .A0(\d0<8> ), .A1(n37), .B0(\d1<8> ), .B1(n39), .Y(n5) );
  OAI2BB1X1 U54 ( .A0N(\d2<10> ), .A1N(n41), .B0(n34), .Y(\y<10> ) );
  OAI2BB1X1 U55 ( .A0N(\d2<11> ), .A1N(n41), .B0(n33), .Y(\y<11> ) );
  OAI2BB1X1 U56 ( .A0N(\d2<12> ), .A1N(n41), .B0(n32), .Y(\y<12> ) );
  OAI2BB1X1 U57 ( .A0N(\d2<13> ), .A1N(n41), .B0(n31), .Y(\y<13> ) );
  OAI2BB1X1 U58 ( .A0N(\d2<14> ), .A1N(n41), .B0(n30), .Y(\y<14> ) );
  OAI2BB1X1 U59 ( .A0N(\d2<15> ), .A1N(n41), .B0(n29), .Y(\y<15> ) );
  OAI2BB1X1 U60 ( .A0N(\d2<16> ), .A1N(n41), .B0(n28), .Y(\y<16> ) );
  OAI2BB1X1 U61 ( .A0N(\d2<17> ), .A1N(n41), .B0(n27), .Y(\y<17> ) );
  OAI2BB1X1 U62 ( .A0N(\d2<18> ), .A1N(n41), .B0(n26), .Y(\y<18> ) );
  OAI2BB1X1 U63 ( .A0N(\d2<19> ), .A1N(n41), .B0(n25), .Y(\y<19> ) );
  OAI2BB1X1 U64 ( .A0N(\d2<20> ), .A1N(n41), .B0(n23), .Y(\y<20> ) );
  OAI2BB1X1 U65 ( .A0N(\d2<21> ), .A1N(n41), .B0(n22), .Y(\y<21> ) );
  OAI2BB1X1 U66 ( .A0N(\d2<22> ), .A1N(n41), .B0(n21), .Y(\y<22> ) );
  OAI2BB1X1 U67 ( .A0N(\d2<23> ), .A1N(n41), .B0(n20), .Y(\y<23> ) );
  OAI2BB1X1 U68 ( .A0N(\d2<24> ), .A1N(n41), .B0(n19), .Y(\y<24> ) );
  OAI2BB1X1 U69 ( .A0N(\d2<25> ), .A1N(n41), .B0(n18), .Y(\y<25> ) );
  OAI2BB1X1 U70 ( .A0N(\d2<26> ), .A1N(n41), .B0(n17), .Y(\y<26> ) );
  OAI2BB1X1 U71 ( .A0N(\d2<27> ), .A1N(n41), .B0(n16), .Y(\y<27> ) );
  OAI2BB1X1 U72 ( .A0N(\d2<28> ), .A1N(n41), .B0(n15), .Y(\y<28> ) );
  OAI2BB1X1 U73 ( .A0N(\d2<29> ), .A1N(n41), .B0(n14), .Y(\y<29> ) );
  OAI2BB1X1 U74 ( .A0N(\d2<30> ), .A1N(n41), .B0(n12), .Y(\y<30> ) );
endmodule


module mux3_WIDTH32_2 ( .d0({\d0<31> , \d0<30> , \d0<29> , \d0<28> , \d0<27> , 
        \d0<26> , \d0<25> , \d0<24> , \d0<23> , \d0<22> , \d0<21> , \d0<20> , 
        \d0<19> , \d0<18> , \d0<17> , \d0<16> , \d0<15> , \d0<14> , \d0<13> , 
        \d0<12> , \d0<11> , \d0<10> , \d0<9> , \d0<8> , \d0<7> , \d0<6> , 
        \d0<5> , \d0<4> , \d0<3> , \d0<2> , \d0<1> , \d0<0> }), .d1({\d1<31> , 
        \d1<30> , \d1<29> , \d1<28> , \d1<27> , \d1<26> , \d1<25> , \d1<24> , 
        \d1<23> , \d1<22> , \d1<21> , \d1<20> , \d1<19> , \d1<18> , \d1<17> , 
        \d1<16> , \d1<15> , \d1<14> , \d1<13> , \d1<12> , \d1<11> , \d1<10> , 
        \d1<9> , \d1<8> , \d1<7> , \d1<6> , \d1<5> , \d1<4> , \d1<3> , \d1<2> , 
        \d1<1> , \d1<0> }), .d2({\d2<31> , \d2<30> , \d2<29> , \d2<28> , 
        \d2<27> , \d2<26> , \d2<25> , \d2<24> , \d2<23> , \d2<22> , \d2<21> , 
        \d2<20> , \d2<19> , \d2<18> , \d2<17> , \d2<16> , \d2<15> , \d2<14> , 
        \d2<13> , \d2<12> , \d2<11> , \d2<10> , \d2<9> , \d2<8> , \d2<7> , 
        \d2<6> , \d2<5> , \d2<4> , \d2<3> , \d2<2> , \d2<1> , \d2<0> }), .s({
        \s<1> , \s<0> }), .y({\y<31> , \y<30> , \y<29> , \y<28> , \y<27> , 
        \y<26> , \y<25> , \y<24> , \y<23> , \y<22> , \y<21> , \y<20> , \y<19> , 
        \y<18> , \y<17> , \y<16> , \y<15> , \y<14> , \y<13> , \y<12> , \y<11> , 
        \y<10> , \y<9> , \y<8> , \y<7> , \y<6> , \y<5> , \y<4> , \y<3> , 
        \y<2> , \y<1> , \y<0> }) );
  input \d0<31> , \d0<30> , \d0<29> , \d0<28> , \d0<27> , \d0<26> , \d0<25> ,
         \d0<24> , \d0<23> , \d0<22> , \d0<21> , \d0<20> , \d0<19> , \d0<18> ,
         \d0<17> , \d0<16> , \d0<15> , \d0<14> , \d0<13> , \d0<12> , \d0<11> ,
         \d0<10> , \d0<9> , \d0<8> , \d0<7> , \d0<6> , \d0<5> , \d0<4> ,
         \d0<3> , \d0<2> , \d0<1> , \d0<0> , \d1<31> , \d1<30> , \d1<29> ,
         \d1<28> , \d1<27> , \d1<26> , \d1<25> , \d1<24> , \d1<23> , \d1<22> ,
         \d1<21> , \d1<20> , \d1<19> , \d1<18> , \d1<17> , \d1<16> , \d1<15> ,
         \d1<14> , \d1<13> , \d1<12> , \d1<11> , \d1<10> , \d1<9> , \d1<8> ,
         \d1<7> , \d1<6> , \d1<5> , \d1<4> , \d1<3> , \d1<2> , \d1<1> ,
         \d1<0> , \d2<31> , \d2<30> , \d2<29> , \d2<28> , \d2<27> , \d2<26> ,
         \d2<25> , \d2<24> , \d2<23> , \d2<22> , \d2<21> , \d2<20> , \d2<19> ,
         \d2<18> , \d2<17> , \d2<16> , \d2<15> , \d2<14> , \d2<13> , \d2<12> ,
         \d2<11> , \d2<10> , \d2<9> , \d2<8> , \d2<7> , \d2<6> , \d2<5> ,
         \d2<4> , \d2<3> , \d2<2> , \d2<1> , \d2<0> , \s<1> , \s<0> ;
  output \y<31> , \y<30> , \y<29> , \y<28> , \y<27> , \y<26> , \y<25> ,
         \y<24> , \y<23> , \y<22> , \y<21> , \y<20> , \y<19> , \y<18> ,
         \y<17> , \y<16> , \y<15> , \y<14> , \y<13> , \y<12> , \y<11> ,
         \y<10> , \y<9> , \y<8> , \y<7> , \y<6> , \y<5> , \y<4> , \y<3> ,
         \y<2> , \y<1> , \y<0> ;
  wire   n1, n3, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61,
         n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75,
         n76;

  INVX12 U1 ( .A(n36), .Y(n1) );
  INVX12 U2 ( .A(n36), .Y(n3) );
  OR2X4 U3 ( .A(\s<0> ), .B(n40), .Y(n36) );
  INVXL U4 ( .A(n75), .Y(n38) );
  OAI2BB1X1 U5 ( .A0N(\d2<1> ), .A1N(n40), .B0(n55), .Y(\y<1> ) );
  AOI22X4 U6 ( .A0(\d0<1> ), .A1(n3), .B0(\d1<1> ), .B1(n75), .Y(n55) );
  CLKINVX3 U7 ( .A(\s<1> ), .Y(n43) );
  INVX16 U8 ( .A(n43), .Y(n40) );
  INVX16 U9 ( .A(n38), .Y(n37) );
  INVX12 U10 ( .A(n36), .Y(n39) );
  OAI2BB1X2 U11 ( .A0N(\d2<2> ), .A1N(n40), .B0(n66), .Y(\y<2> ) );
  AOI22X1 U12 ( .A0(\d0<2> ), .A1(n39), .B0(\d1<2> ), .B1(n75), .Y(n66) );
  OAI2BB1X1 U13 ( .A0N(\d2<3> ), .A1N(n40), .B0(n69), .Y(\y<3> ) );
  OAI2BB1X1 U14 ( .A0N(\d2<4> ), .A1N(n40), .B0(n70), .Y(\y<4> ) );
  AOI22X2 U15 ( .A0(\d0<0> ), .A1(n1), .B0(\d1<0> ), .B1(n75), .Y(n44) );
  INVXL U16 ( .A(n40), .Y(n42) );
  AOI22XL U17 ( .A0(\d0<4> ), .A1(n39), .B0(\d1<4> ), .B1(n75), .Y(n70) );
  AOI22XL U18 ( .A0(\d0<16> ), .A1(n3), .B0(\d1<16> ), .B1(n37), .Y(n51) );
  AOI22XL U19 ( .A0(\d0<15> ), .A1(n39), .B0(\d1<15> ), .B1(n37), .Y(n50) );
  AOI22XL U20 ( .A0(\d0<14> ), .A1(n3), .B0(\d1<14> ), .B1(n37), .Y(n49) );
  AOI22XL U21 ( .A0(\d0<20> ), .A1(n39), .B0(\d1<20> ), .B1(n37), .Y(n56) );
  AOI22XL U22 ( .A0(\d0<19> ), .A1(n3), .B0(\d1<19> ), .B1(n37), .Y(n54) );
  AOI22XL U23 ( .A0(\d0<18> ), .A1(n39), .B0(\d1<18> ), .B1(n37), .Y(n53) );
  AOI22XL U24 ( .A0(\d0<17> ), .A1(n39), .B0(\d1<17> ), .B1(n37), .Y(n52) );
  AOI22XL U25 ( .A0(\d0<24> ), .A1(n3), .B0(\d1<24> ), .B1(n37), .Y(n60) );
  AOI22XL U26 ( .A0(\d0<23> ), .A1(n39), .B0(\d1<23> ), .B1(n37), .Y(n59) );
  AOI22XL U27 ( .A0(\d0<22> ), .A1(n1), .B0(\d1<22> ), .B1(n37), .Y(n58) );
  AOI22XL U28 ( .A0(\d0<21> ), .A1(n3), .B0(\d1<21> ), .B1(n37), .Y(n57) );
  AOI22XL U29 ( .A0(\d0<26> ), .A1(n1), .B0(\d1<26> ), .B1(n37), .Y(n62) );
  AOI22XL U30 ( .A0(\d0<25> ), .A1(n39), .B0(\d1<25> ), .B1(n37), .Y(n61) );
  AOI22XL U31 ( .A0(\d0<30> ), .A1(n3), .B0(\d1<30> ), .B1(n37), .Y(n67) );
  NOR2BX4 U32 ( .AN(\s<0> ), .B(n40), .Y(n75) );
  OAI2BB1X4 U33 ( .A0N(\d2<0> ), .A1N(n40), .B0(n44), .Y(\y<0> ) );
  CLKINVX3 U34 ( .A(n42), .Y(n41) );
  AOI22X1 U35 ( .A0(\d0<3> ), .A1(n39), .B0(\d1<3> ), .B1(n75), .Y(n69) );
  OAI2BB1X1 U36 ( .A0N(\d2<5> ), .A1N(n40), .B0(n71), .Y(\y<5> ) );
  AOI22X1 U37 ( .A0(\d0<5> ), .A1(n39), .B0(\d1<5> ), .B1(n37), .Y(n71) );
  OAI2BB1X1 U38 ( .A0N(\d2<6> ), .A1N(n40), .B0(n72), .Y(\y<6> ) );
  AOI22X1 U39 ( .A0(\d0<6> ), .A1(n39), .B0(\d1<6> ), .B1(n37), .Y(n72) );
  OAI2BB1X1 U40 ( .A0N(\d2<7> ), .A1N(n40), .B0(n73), .Y(\y<7> ) );
  AOI22X1 U41 ( .A0(\d0<7> ), .A1(n39), .B0(\d1<7> ), .B1(n37), .Y(n73) );
  OAI2BB1X1 U42 ( .A0N(\d2<8> ), .A1N(n40), .B0(n74), .Y(\y<8> ) );
  AOI22X1 U43 ( .A0(\d0<8> ), .A1(n39), .B0(\d1<8> ), .B1(n37), .Y(n74) );
  OAI2BB1X1 U44 ( .A0N(n40), .A1N(\d2<9> ), .B0(n76), .Y(\y<9> ) );
  AOI22X1 U45 ( .A0(\d0<9> ), .A1(n39), .B0(\d1<9> ), .B1(n37), .Y(n76) );
  OAI2BB1X1 U46 ( .A0N(\d2<10> ), .A1N(n40), .B0(n45), .Y(\y<10> ) );
  AOI22X1 U47 ( .A0(\d0<10> ), .A1(n39), .B0(\d1<10> ), .B1(n37), .Y(n45) );
  OAI2BB1X1 U48 ( .A0N(\d2<11> ), .A1N(n40), .B0(n46), .Y(\y<11> ) );
  AOI22X1 U49 ( .A0(\d0<11> ), .A1(n39), .B0(\d1<11> ), .B1(n37), .Y(n46) );
  OAI2BB1X1 U50 ( .A0N(\d2<12> ), .A1N(n40), .B0(n47), .Y(\y<12> ) );
  AOI22X1 U51 ( .A0(\d0<12> ), .A1(n3), .B0(\d1<12> ), .B1(n37), .Y(n47) );
  OAI2BB1X1 U52 ( .A0N(\d2<13> ), .A1N(n41), .B0(n48), .Y(\y<13> ) );
  AOI22X1 U53 ( .A0(\d0<13> ), .A1(n39), .B0(\d1<13> ), .B1(n37), .Y(n48) );
  OAI2BB1X1 U54 ( .A0N(\d2<14> ), .A1N(n41), .B0(n49), .Y(\y<14> ) );
  OAI2BB1X1 U55 ( .A0N(\d2<15> ), .A1N(n41), .B0(n50), .Y(\y<15> ) );
  OAI2BB1X1 U56 ( .A0N(\d2<16> ), .A1N(n41), .B0(n51), .Y(\y<16> ) );
  OAI2BB1X1 U57 ( .A0N(\d2<17> ), .A1N(n41), .B0(n52), .Y(\y<17> ) );
  OAI2BB1X1 U58 ( .A0N(\d2<18> ), .A1N(n41), .B0(n53), .Y(\y<18> ) );
  OAI2BB1X1 U59 ( .A0N(\d2<19> ), .A1N(n41), .B0(n54), .Y(\y<19> ) );
  OAI2BB1X1 U60 ( .A0N(\d2<20> ), .A1N(n41), .B0(n56), .Y(\y<20> ) );
  OAI2BB1X1 U61 ( .A0N(\d2<21> ), .A1N(n41), .B0(n57), .Y(\y<21> ) );
  OAI2BB1X1 U62 ( .A0N(\d2<22> ), .A1N(n41), .B0(n58), .Y(\y<22> ) );
  OAI2BB1X1 U63 ( .A0N(\d2<25> ), .A1N(n41), .B0(n61), .Y(\y<25> ) );
  OAI2BB1X1 U64 ( .A0N(\d2<23> ), .A1N(n41), .B0(n59), .Y(\y<23> ) );
  OAI2BB1X1 U65 ( .A0N(\d2<24> ), .A1N(n41), .B0(n60), .Y(\y<24> ) );
  OAI2BB1X1 U66 ( .A0N(\d2<26> ), .A1N(n41), .B0(n62), .Y(\y<26> ) );
  OAI2BB1X1 U67 ( .A0N(\d2<27> ), .A1N(n40), .B0(n63), .Y(\y<27> ) );
  AOI22X1 U68 ( .A0(\d0<27> ), .A1(n3), .B0(\d1<27> ), .B1(n37), .Y(n63) );
  OAI2BB1X1 U69 ( .A0N(\d2<28> ), .A1N(n40), .B0(n64), .Y(\y<28> ) );
  AOI22X1 U70 ( .A0(\d0<28> ), .A1(n39), .B0(\d1<28> ), .B1(n37), .Y(n64) );
  OAI2BB1X1 U71 ( .A0N(\d2<31> ), .A1N(n40), .B0(n68), .Y(\y<31> ) );
  AOI22X1 U72 ( .A0(\d0<31> ), .A1(n39), .B0(\d1<31> ), .B1(n37), .Y(n68) );
  OAI2BB1X1 U73 ( .A0N(\d2<29> ), .A1N(n40), .B0(n65), .Y(\y<29> ) );
  AOI22X1 U74 ( .A0(\d0<29> ), .A1(n1), .B0(\d1<29> ), .B1(n37), .Y(n65) );
  OAI2BB1X1 U75 ( .A0N(\d2<30> ), .A1N(n41), .B0(n67), .Y(\y<30> ) );
endmodule


module mux3_WIDTH32_1 ( .d0({\d0<31> , \d0<30> , \d0<29> , \d0<28> , \d0<27> , 
        \d0<26> , \d0<25> , \d0<24> , \d0<23> , \d0<22> , \d0<21> , \d0<20> , 
        \d0<19> , \d0<18> , \d0<17> , \d0<16> , \d0<15> , \d0<14> , \d0<13> , 
        \d0<12> , \d0<11> , \d0<10> , \d0<9> , \d0<8> , \d0<7> , \d0<6> , 
        \d0<5> , \d0<4> , \d0<3> , \d0<2> , \d0<1> , \d0<0> }), .d1({\d1<31> , 
        \d1<30> , \d1<29> , \d1<28> , \d1<27> , \d1<26> , \d1<25> , \d1<24> , 
        \d1<23> , \d1<22> , \d1<21> , \d1<20> , \d1<19> , \d1<18> , \d1<17> , 
        \d1<16> , \d1<15> , \d1<14> , \d1<13> , \d1<12> , \d1<11> , \d1<10> , 
        \d1<9> , \d1<8> , \d1<7> , \d1<6> , \d1<5> , \d1<4> , \d1<3> , \d1<2> , 
        \d1<1> , \d1<0> }), .d2({\d2<31> , \d2<30> , \d2<29> , \d2<28> , 
        \d2<27> , \d2<26> , \d2<25> , \d2<24> , \d2<23> , \d2<22> , \d2<21> , 
        \d2<20> , \d2<19> , \d2<18> , \d2<17> , \d2<16> , \d2<15> , \d2<14> , 
        \d2<13> , \d2<12> , \d2<11> , \d2<10> , \d2<9> , \d2<8> , \d2<7> , 
        \d2<6> , \d2<5> , \d2<4> , \d2<3> , \d2<2> , \d2<1> , \d2<0> }), .s({
        \s<1> , \s<0> }), .y({\y<31> , \y<30> , \y<29> , \y<28> , \y<27> , 
        \y<26> , \y<25> , \y<24> , \y<23> , \y<22> , \y<21> , \y<20> , \y<19> , 
        \y<18> , \y<17> , \y<16> , \y<15> , \y<14> , \y<13> , \y<12> , \y<11> , 
        \y<10> , \y<9> , \y<8> , \y<7> , \y<6> , \y<5> , \y<4> , \y<3> , 
        \y<2> , \y<1> , \y<0> }) );
  input \d0<31> , \d0<30> , \d0<29> , \d0<28> , \d0<27> , \d0<26> , \d0<25> ,
         \d0<24> , \d0<23> , \d0<22> , \d0<21> , \d0<20> , \d0<19> , \d0<18> ,
         \d0<17> , \d0<16> , \d0<15> , \d0<14> , \d0<13> , \d0<12> , \d0<11> ,
         \d0<10> , \d0<9> , \d0<8> , \d0<7> , \d0<6> , \d0<5> , \d0<4> ,
         \d0<3> , \d0<2> , \d0<1> , \d0<0> , \d1<31> , \d1<30> , \d1<29> ,
         \d1<28> , \d1<27> , \d1<26> , \d1<25> , \d1<24> , \d1<23> , \d1<22> ,
         \d1<21> , \d1<20> , \d1<19> , \d1<18> , \d1<17> , \d1<16> , \d1<15> ,
         \d1<14> , \d1<13> , \d1<12> , \d1<11> , \d1<10> , \d1<9> , \d1<8> ,
         \d1<7> , \d1<6> , \d1<5> , \d1<4> , \d1<3> , \d1<2> , \d1<1> ,
         \d1<0> , \d2<31> , \d2<30> , \d2<29> , \d2<28> , \d2<27> , \d2<26> ,
         \d2<25> , \d2<24> , \d2<23> , \d2<22> , \d2<21> , \d2<20> , \d2<19> ,
         \d2<18> , \d2<17> , \d2<16> , \d2<15> , \d2<14> , \d2<13> , \d2<12> ,
         \d2<11> , \d2<10> , \d2<9> , \d2<8> , \d2<7> , \d2<6> , \d2<5> ,
         \d2<4> , \d2<3> , \d2<2> , \d2<1> , \d2<0> , \s<1> , \s<0> ;
  output \y<31> , \y<30> , \y<29> , \y<28> , \y<27> , \y<26> , \y<25> ,
         \y<24> , \y<23> , \y<22> , \y<21> , \y<20> , \y<19> , \y<18> ,
         \y<17> , \y<16> , \y<15> , \y<14> , \y<13> , \y<12> , \y<11> ,
         \y<10> , \y<9> , \y<8> , \y<7> , \y<6> , \y<5> , \y<4> , \y<3> ,
         \y<2> , \y<1> , \y<0> ;
  wire   n1, n3, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61,
         n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75;

  OAI2BB1X4 U1 ( .A0N(\d2<26> ), .A1N(n41), .B0(n61), .Y(\y<26> ) );
  OAI2BB1X1 U2 ( .A0N(\d2<30> ), .A1N(n41), .B0(n66), .Y(\y<30> ) );
  OAI2BB1X4 U3 ( .A0N(\d2<31> ), .A1N(n40), .B0(n67), .Y(\y<31> ) );
  OAI2BB1X4 U4 ( .A0N(\d2<27> ), .A1N(n40), .B0(n62), .Y(\y<27> ) );
  OAI2BB1X1 U5 ( .A0N(\d2<17> ), .A1N(n41), .B0(n51), .Y(\y<17> ) );
  OAI2BB1X1 U6 ( .A0N(\d2<18> ), .A1N(n41), .B0(n52), .Y(\y<18> ) );
  OAI2BB1X1 U7 ( .A0N(\d2<19> ), .A1N(n41), .B0(n53), .Y(\y<19> ) );
  OAI2BB1X1 U8 ( .A0N(\d2<20> ), .A1N(n41), .B0(n55), .Y(\y<20> ) );
  OAI2BB1X1 U9 ( .A0N(\d2<21> ), .A1N(n41), .B0(n56), .Y(\y<21> ) );
  OAI2BB1X1 U10 ( .A0N(\d2<22> ), .A1N(n41), .B0(n57), .Y(\y<22> ) );
  OAI2BB1X1 U11 ( .A0N(\d2<24> ), .A1N(n41), .B0(n59), .Y(\y<24> ) );
  OAI2BB1X1 U12 ( .A0N(\d2<25> ), .A1N(n41), .B0(n60), .Y(\y<25> ) );
  OAI2BB1X2 U13 ( .A0N(\d2<28> ), .A1N(n40), .B0(n63), .Y(\y<28> ) );
  OAI2BB1X2 U14 ( .A0N(\d2<29> ), .A1N(n40), .B0(n64), .Y(\y<29> ) );
  OAI2BB1X1 U15 ( .A0N(\d2<10> ), .A1N(n41), .B0(n44), .Y(\y<10> ) );
  OR2X2 U16 ( .A(\s<0> ), .B(n40), .Y(n1) );
  OAI2BB1X1 U17 ( .A0N(\d2<16> ), .A1N(n41), .B0(n50), .Y(\y<16> ) );
  OAI2BB1X1 U18 ( .A0N(\d2<11> ), .A1N(n41), .B0(n45), .Y(\y<11> ) );
  OAI2BB1X4 U19 ( .A0N(\d2<23> ), .A1N(n41), .B0(n58), .Y(\y<23> ) );
  OAI2BB1X4 U20 ( .A0N(\d2<15> ), .A1N(n41), .B0(n49), .Y(\y<15> ) );
  OAI2BB1X4 U21 ( .A0N(\d2<14> ), .A1N(n41), .B0(n48), .Y(\y<14> ) );
  OAI2BB1X4 U22 ( .A0N(\d2<13> ), .A1N(n41), .B0(n47), .Y(\y<13> ) );
  OAI2BB1X4 U23 ( .A0N(\d2<12> ), .A1N(n41), .B0(n46), .Y(\y<12> ) );
  OAI2BB1X1 U24 ( .A0N(\d2<8> ), .A1N(n40), .B0(n73), .Y(\y<8> ) );
  OAI2BB1X1 U25 ( .A0N(n40), .A1N(\d2<9> ), .B0(n75), .Y(\y<9> ) );
  OAI2BB1X1 U26 ( .A0N(\d2<7> ), .A1N(n40), .B0(n72), .Y(\y<7> ) );
  OAI2BB1X1 U27 ( .A0N(\d2<6> ), .A1N(n40), .B0(n71), .Y(\y<6> ) );
  OAI2BB1X1 U28 ( .A0N(\d2<5> ), .A1N(n40), .B0(n70), .Y(\y<5> ) );
  OAI2BB1X1 U29 ( .A0N(\d2<0> ), .A1N(n40), .B0(n43), .Y(\y<0> ) );
  OAI2BB1X1 U30 ( .A0N(\d2<2> ), .A1N(n40), .B0(n65), .Y(\y<2> ) );
  OAI2BB1X1 U31 ( .A0N(\d2<1> ), .A1N(n41), .B0(n54), .Y(\y<1> ) );
  OAI2BB1X1 U32 ( .A0N(\d2<4> ), .A1N(n40), .B0(n69), .Y(\y<4> ) );
  OAI2BB1X1 U33 ( .A0N(\d2<3> ), .A1N(n40), .B0(n68), .Y(\y<3> ) );
  AOI22XL U34 ( .A0(\d0<0> ), .A1(n39), .B0(\d1<0> ), .B1(n3), .Y(n43) );
  AOI22XL U35 ( .A0(\d0<2> ), .A1(n38), .B0(\d1<2> ), .B1(n36), .Y(n65) );
  AOI22XL U36 ( .A0(\d0<1> ), .A1(n39), .B0(\d1<1> ), .B1(n3), .Y(n54) );
  CLKINVX3 U37 ( .A(n42), .Y(n41) );
  CLKINVX3 U38 ( .A(n42), .Y(n40) );
  INVX1 U39 ( .A(\s<1> ), .Y(n42) );
  CLKINVX3 U40 ( .A(n1), .Y(n38) );
  CLKINVX3 U41 ( .A(n37), .Y(n36) );
  CLKINVX3 U42 ( .A(n1), .Y(n39) );
  CLKINVX3 U43 ( .A(n37), .Y(n3) );
  INVX1 U44 ( .A(n74), .Y(n37) );
  NOR2BX1 U45 ( .AN(\s<0> ), .B(n40), .Y(n74) );
  AOI22X1 U46 ( .A0(\d0<31> ), .A1(n39), .B0(\d1<31> ), .B1(n36), .Y(n67) );
  AOI22X1 U47 ( .A0(\d0<26> ), .A1(n38), .B0(\d1<26> ), .B1(n36), .Y(n61) );
  AOI22X1 U48 ( .A0(\d0<27> ), .A1(n38), .B0(\d1<27> ), .B1(n36), .Y(n62) );
  AOI22X1 U49 ( .A0(\d0<28> ), .A1(n38), .B0(\d1<28> ), .B1(n36), .Y(n63) );
  AOI22X1 U50 ( .A0(\d0<29> ), .A1(n38), .B0(\d1<29> ), .B1(n36), .Y(n64) );
  AOI22X1 U51 ( .A0(\d0<30> ), .A1(n38), .B0(\d1<30> ), .B1(n36), .Y(n66) );
  AOI22X1 U52 ( .A0(\d0<21> ), .A1(n38), .B0(\d1<21> ), .B1(n36), .Y(n56) );
  AOI22X1 U53 ( .A0(\d0<22> ), .A1(n38), .B0(\d1<22> ), .B1(n36), .Y(n57) );
  AOI22X1 U54 ( .A0(\d0<23> ), .A1(n38), .B0(\d1<23> ), .B1(n36), .Y(n58) );
  AOI22X1 U55 ( .A0(\d0<24> ), .A1(n38), .B0(\d1<24> ), .B1(n36), .Y(n59) );
  AOI22X1 U56 ( .A0(\d0<25> ), .A1(n38), .B0(\d1<25> ), .B1(n36), .Y(n60) );
  AOI22X1 U57 ( .A0(\d0<16> ), .A1(n39), .B0(\d1<16> ), .B1(n3), .Y(n50) );
  AOI22X1 U58 ( .A0(\d0<17> ), .A1(n39), .B0(\d1<17> ), .B1(n3), .Y(n51) );
  AOI22X1 U59 ( .A0(\d0<18> ), .A1(n38), .B0(\d1<18> ), .B1(n3), .Y(n52) );
  AOI22X1 U60 ( .A0(\d0<19> ), .A1(n39), .B0(\d1<19> ), .B1(n3), .Y(n53) );
  AOI22X1 U61 ( .A0(\d0<20> ), .A1(n38), .B0(\d1<20> ), .B1(n36), .Y(n55) );
  AOI22X1 U62 ( .A0(\d0<10> ), .A1(n38), .B0(\d1<10> ), .B1(n3), .Y(n44) );
  AOI22X1 U63 ( .A0(\d0<11> ), .A1(n39), .B0(\d1<11> ), .B1(n3), .Y(n45) );
  AOI22X1 U64 ( .A0(\d0<12> ), .A1(n39), .B0(\d1<12> ), .B1(n3), .Y(n46) );
  AOI22X1 U65 ( .A0(\d0<13> ), .A1(n38), .B0(\d1<13> ), .B1(n3), .Y(n47) );
  AOI22X1 U66 ( .A0(\d0<14> ), .A1(n39), .B0(\d1<14> ), .B1(n3), .Y(n48) );
  AOI22X1 U67 ( .A0(\d0<15> ), .A1(n38), .B0(\d1<15> ), .B1(n3), .Y(n49) );
  AOI22X1 U68 ( .A0(\d0<9> ), .A1(n39), .B0(\d1<9> ), .B1(n3), .Y(n75) );
  AOI22X1 U69 ( .A0(\d0<5> ), .A1(n39), .B0(\d1<5> ), .B1(n3), .Y(n70) );
  AOI22X1 U70 ( .A0(\d0<6> ), .A1(n39), .B0(\d1<6> ), .B1(n36), .Y(n71) );
  AOI22X1 U71 ( .A0(\d0<7> ), .A1(n39), .B0(\d1<7> ), .B1(n3), .Y(n72) );
  AOI22X1 U72 ( .A0(\d0<8> ), .A1(n39), .B0(\d1<8> ), .B1(n36), .Y(n73) );
  AOI22X1 U73 ( .A0(\d0<3> ), .A1(n39), .B0(\d1<3> ), .B1(n3), .Y(n68) );
  AOI22X1 U74 ( .A0(\d0<4> ), .A1(n39), .B0(\d1<4> ), .B1(n36), .Y(n69) );
endmodule


module regfile ( clk, we3, .ra1({\ra1<3> , \ra1<2> , \ra1<1> , \ra1<0> }), 
    .ra2({\ra2<3> , \ra2<2> , \ra2<1> , \ra2<0> }), .wa3({\wa3<3> , \wa3<2> , 
        \wa3<1> , \wa3<0> }), .wd3({\wd3<31> , \wd3<30> , \wd3<29> , \wd3<28> , 
        \wd3<27> , \wd3<26> , \wd3<25> , \wd3<24> , \wd3<23> , \wd3<22> , 
        \wd3<21> , \wd3<20> , \wd3<19> , \wd3<18> , \wd3<17> , \wd3<16> , 
        \wd3<15> , \wd3<14> , \wd3<13> , \wd3<12> , \wd3<11> , \wd3<10> , 
        \wd3<9> , \wd3<8> , \wd3<7> , \wd3<6> , \wd3<5> , \wd3<4> , \wd3<3> , 
        \wd3<2> , \wd3<1> , \wd3<0> }), .r15({\r15<31> , \r15<30> , \r15<29> , 
        \r15<28> , \r15<27> , \r15<26> , \r15<25> , \r15<24> , \r15<23> , 
        \r15<22> , \r15<21> , \r15<20> , \r15<19> , \r15<18> , \r15<17> , 
        \r15<16> , \r15<15> , \r15<14> , \r15<13> , \r15<12> , \r15<11> , 
        \r15<10> , \r15<9> , \r15<8> , \r15<7> , \r15<6> , \r15<5> , \r15<4> , 
        \r15<3> , \r15<2> , \r15<1> , \r15<0> }), .rd1({\rd1<31> , \rd1<30> , 
        \rd1<29> , \rd1<28> , \rd1<27> , \rd1<26> , \rd1<25> , \rd1<24> , 
        \rd1<23> , \rd1<22> , \rd1<21> , \rd1<20> , \rd1<19> , \rd1<18> , 
        \rd1<17> , \rd1<16> , \rd1<15> , \rd1<14> , \rd1<13> , \rd1<12> , 
        \rd1<11> , \rd1<10> , \rd1<9> , \rd1<8> , \rd1<7> , \rd1<6> , \rd1<5> , 
        \rd1<4> , \rd1<3> , \rd1<2> , \rd1<1> , \rd1<0> }), .rd2({\rd2<31> , 
        \rd2<30> , \rd2<29> , \rd2<28> , \rd2<27> , \rd2<26> , \rd2<25> , 
        \rd2<24> , \rd2<23> , \rd2<22> , \rd2<21> , \rd2<20> , \rd2<19> , 
        \rd2<18> , \rd2<17> , \rd2<16> , \rd2<15> , \rd2<14> , \rd2<13> , 
        \rd2<12> , \rd2<11> , \rd2<10> , \rd2<9> , \rd2<8> , \rd2<7> , 
        \rd2<6> , \rd2<5> , \rd2<4> , \rd2<3> , \rd2<2> , \rd2<1> , \rd2<0> })
 );
  input clk, we3, \ra1<3> , \ra1<2> , \ra1<1> , \ra1<0> , \ra2<3> , \ra2<2> ,
         \ra2<1> , \ra2<0> , \wa3<3> , \wa3<2> , \wa3<1> , \wa3<0> , \wd3<31> ,
         \wd3<30> , \wd3<29> , \wd3<28> , \wd3<27> , \wd3<26> , \wd3<25> ,
         \wd3<24> , \wd3<23> , \wd3<22> , \wd3<21> , \wd3<20> , \wd3<19> ,
         \wd3<18> , \wd3<17> , \wd3<16> , \wd3<15> , \wd3<14> , \wd3<13> ,
         \wd3<12> , \wd3<11> , \wd3<10> , \wd3<9> , \wd3<8> , \wd3<7> ,
         \wd3<6> , \wd3<5> , \wd3<4> , \wd3<3> , \wd3<2> , \wd3<1> , \wd3<0> ,
         \r15<31> , \r15<30> , \r15<29> , \r15<28> , \r15<27> , \r15<26> ,
         \r15<25> , \r15<24> , \r15<23> , \r15<22> , \r15<21> , \r15<20> ,
         \r15<19> , \r15<18> , \r15<17> , \r15<16> , \r15<15> , \r15<14> ,
         \r15<13> , \r15<12> , \r15<11> , \r15<10> , \r15<9> , \r15<8> ,
         \r15<7> , \r15<6> , \r15<5> , \r15<4> , \r15<3> , \r15<2> , \r15<1> ,
         \r15<0> ;
  output \rd1<31> , \rd1<30> , \rd1<29> , \rd1<28> , \rd1<27> , \rd1<26> ,
         \rd1<25> , \rd1<24> , \rd1<23> , \rd1<22> , \rd1<21> , \rd1<20> ,
         \rd1<19> , \rd1<18> , \rd1<17> , \rd1<16> , \rd1<15> , \rd1<14> ,
         \rd1<13> , \rd1<12> , \rd1<11> , \rd1<10> , \rd1<9> , \rd1<8> ,
         \rd1<7> , \rd1<6> , \rd1<5> , \rd1<4> , \rd1<3> , \rd1<2> , \rd1<1> ,
         \rd1<0> , \rd2<31> , \rd2<30> , \rd2<29> , \rd2<28> , \rd2<27> ,
         \rd2<26> , \rd2<25> , \rd2<24> , \rd2<23> , \rd2<22> , \rd2<21> ,
         \rd2<20> , \rd2<19> , \rd2<18> , \rd2<17> , \rd2<16> , \rd2<15> ,
         \rd2<14> , \rd2<13> , \rd2<12> , \rd2<11> , \rd2<10> , \rd2<9> ,
         \rd2<8> , \rd2<7> , \rd2<6> , \rd2<5> , \rd2<4> , \rd2<3> , \rd2<2> ,
         \rd2<1> , \rd2<0> ;
  wire   N12, N13, N14, N15, N16, N17, N18, N19, \rf<14><31> , \rf<14><30> ,
         \rf<14><29> , \rf<14><28> , \rf<14><27> , \rf<14><26> , \rf<14><25> ,
         \rf<14><24> , \rf<14><23> , \rf<14><22> , \rf<14><21> , \rf<14><20> ,
         \rf<14><19> , \rf<14><18> , \rf<14><17> , \rf<14><16> , \rf<14><15> ,
         \rf<14><14> , \rf<14><13> , \rf<14><12> , \rf<14><11> , \rf<14><10> ,
         \rf<14><9> , \rf<14><8> , \rf<14><7> , \rf<14><6> , \rf<14><5> ,
         \rf<14><4> , \rf<14><3> , \rf<14><2> , \rf<14><1> , \rf<14><0> ,
         \rf<13><31> , \rf<13><30> , \rf<13><29> , \rf<13><28> , \rf<13><27> ,
         \rf<13><26> , \rf<13><25> , \rf<13><24> , \rf<13><23> , \rf<13><22> ,
         \rf<13><21> , \rf<13><20> , \rf<13><19> , \rf<13><18> , \rf<13><17> ,
         \rf<13><16> , \rf<13><15> , \rf<13><14> , \rf<13><13> , \rf<13><12> ,
         \rf<13><11> , \rf<13><10> , \rf<13><9> , \rf<13><8> , \rf<13><7> ,
         \rf<13><6> , \rf<13><5> , \rf<13><4> , \rf<13><3> , \rf<13><2> ,
         \rf<13><1> , \rf<13><0> , \rf<12><31> , \rf<12><30> , \rf<12><29> ,
         \rf<12><28> , \rf<12><27> , \rf<12><26> , \rf<12><25> , \rf<12><24> ,
         \rf<12><23> , \rf<12><22> , \rf<12><21> , \rf<12><20> , \rf<12><19> ,
         \rf<12><18> , \rf<12><17> , \rf<12><16> , \rf<12><15> , \rf<12><14> ,
         \rf<12><13> , \rf<12><12> , \rf<12><11> , \rf<12><10> , \rf<12><9> ,
         \rf<12><8> , \rf<12><7> , \rf<12><6> , \rf<12><5> , \rf<12><4> ,
         \rf<12><3> , \rf<12><2> , \rf<12><1> , \rf<12><0> , \rf<11><31> ,
         \rf<11><30> , \rf<11><29> , \rf<11><28> , \rf<11><27> , \rf<11><26> ,
         \rf<11><25> , \rf<11><24> , \rf<11><23> , \rf<11><22> , \rf<11><21> ,
         \rf<11><20> , \rf<11><19> , \rf<11><18> , \rf<11><17> , \rf<11><16> ,
         \rf<11><15> , \rf<11><14> , \rf<11><13> , \rf<11><12> , \rf<11><11> ,
         \rf<11><10> , \rf<11><9> , \rf<11><8> , \rf<11><7> , \rf<11><6> ,
         \rf<11><5> , \rf<11><4> , \rf<11><3> , \rf<11><2> , \rf<11><1> ,
         \rf<11><0> , \rf<10><31> , \rf<10><30> , \rf<10><29> , \rf<10><28> ,
         \rf<10><27> , \rf<10><26> , \rf<10><25> , \rf<10><24> , \rf<10><23> ,
         \rf<10><22> , \rf<10><21> , \rf<10><20> , \rf<10><19> , \rf<10><18> ,
         \rf<10><17> , \rf<10><16> , \rf<10><15> , \rf<10><14> , \rf<10><13> ,
         \rf<10><12> , \rf<10><11> , \rf<10><10> , \rf<10><9> , \rf<10><8> ,
         \rf<10><7> , \rf<10><6> , \rf<10><5> , \rf<10><4> , \rf<10><3> ,
         \rf<10><2> , \rf<10><1> , \rf<10><0> , \rf<9><31> , \rf<9><30> ,
         \rf<9><29> , \rf<9><28> , \rf<9><27> , \rf<9><26> , \rf<9><25> ,
         \rf<9><24> , \rf<9><23> , \rf<9><22> , \rf<9><21> , \rf<9><20> ,
         \rf<9><19> , \rf<9><18> , \rf<9><17> , \rf<9><16> , \rf<9><15> ,
         \rf<9><14> , \rf<9><13> , \rf<9><12> , \rf<9><11> , \rf<9><10> ,
         \rf<9><9> , \rf<9><8> , \rf<9><7> , \rf<9><6> , \rf<9><5> ,
         \rf<9><4> , \rf<9><3> , \rf<9><2> , \rf<9><1> , \rf<9><0> ,
         \rf<8><31> , \rf<8><30> , \rf<8><29> , \rf<8><28> , \rf<8><27> ,
         \rf<8><26> , \rf<8><25> , \rf<8><24> , \rf<8><23> , \rf<8><22> ,
         \rf<8><21> , \rf<8><20> , \rf<8><19> , \rf<8><18> , \rf<8><17> ,
         \rf<8><16> , \rf<8><15> , \rf<8><14> , \rf<8><13> , \rf<8><12> ,
         \rf<8><11> , \rf<8><10> , \rf<8><9> , \rf<8><8> , \rf<8><7> ,
         \rf<8><6> , \rf<8><5> , \rf<8><4> , \rf<8><3> , \rf<8><2> ,
         \rf<8><1> , \rf<8><0> , \rf<7><31> , \rf<7><30> , \rf<7><29> ,
         \rf<7><28> , \rf<7><27> , \rf<7><26> , \rf<7><25> , \rf<7><24> ,
         \rf<7><23> , \rf<7><22> , \rf<7><21> , \rf<7><20> , \rf<7><19> ,
         \rf<7><18> , \rf<7><17> , \rf<7><16> , \rf<7><15> , \rf<7><14> ,
         \rf<7><13> , \rf<7><12> , \rf<7><11> , \rf<7><10> , \rf<7><9> ,
         \rf<7><8> , \rf<7><7> , \rf<7><6> , \rf<7><5> , \rf<7><4> ,
         \rf<7><3> , \rf<7><2> , \rf<7><1> , \rf<7><0> , \rf<6><31> ,
         \rf<6><30> , \rf<6><29> , \rf<6><28> , \rf<6><27> , \rf<6><26> ,
         \rf<6><25> , \rf<6><24> , \rf<6><23> , \rf<6><22> , \rf<6><21> ,
         \rf<6><20> , \rf<6><19> , \rf<6><18> , \rf<6><17> , \rf<6><16> ,
         \rf<6><15> , \rf<6><14> , \rf<6><13> , \rf<6><12> , \rf<6><11> ,
         \rf<6><10> , \rf<6><9> , \rf<6><8> , \rf<6><7> , \rf<6><6> ,
         \rf<6><5> , \rf<6><4> , \rf<6><3> , \rf<6><2> , \rf<6><1> ,
         \rf<6><0> , \rf<5><31> , \rf<5><30> , \rf<5><29> , \rf<5><28> ,
         \rf<5><27> , \rf<5><26> , \rf<5><25> , \rf<5><24> , \rf<5><23> ,
         \rf<5><22> , \rf<5><21> , \rf<5><20> , \rf<5><19> , \rf<5><18> ,
         \rf<5><17> , \rf<5><16> , \rf<5><15> , \rf<5><14> , \rf<5><13> ,
         \rf<5><12> , \rf<5><11> , \rf<5><10> , \rf<5><9> , \rf<5><8> ,
         \rf<5><7> , \rf<5><6> , \rf<5><5> , \rf<5><4> , \rf<5><3> ,
         \rf<5><2> , \rf<5><1> , \rf<5><0> , \rf<4><31> , \rf<4><30> ,
         \rf<4><29> , \rf<4><28> , \rf<4><27> , \rf<4><26> , \rf<4><25> ,
         \rf<4><24> , \rf<4><23> , \rf<4><22> , \rf<4><21> , \rf<4><20> ,
         \rf<4><19> , \rf<4><18> , \rf<4><17> , \rf<4><16> , \rf<4><15> ,
         \rf<4><14> , \rf<4><13> , \rf<4><12> , \rf<4><11> , \rf<4><10> ,
         \rf<4><9> , \rf<4><8> , \rf<4><7> , \rf<4><6> , \rf<4><5> ,
         \rf<4><4> , \rf<4><3> , \rf<4><2> , \rf<4><1> , \rf<4><0> ,
         \rf<3><31> , \rf<3><30> , \rf<3><29> , \rf<3><28> , \rf<3><27> ,
         \rf<3><26> , \rf<3><25> , \rf<3><24> , \rf<3><23> , \rf<3><22> ,
         \rf<3><21> , \rf<3><20> , \rf<3><19> , \rf<3><18> , \rf<3><17> ,
         \rf<3><16> , \rf<3><15> , \rf<3><14> , \rf<3><13> , \rf<3><12> ,
         \rf<3><11> , \rf<3><10> , \rf<3><9> , \rf<3><8> , \rf<3><7> ,
         \rf<3><6> , \rf<3><5> , \rf<3><4> , \rf<3><3> , \rf<3><2> ,
         \rf<3><1> , \rf<3><0> , \rf<2><31> , \rf<2><30> , \rf<2><29> ,
         \rf<2><28> , \rf<2><27> , \rf<2><26> , \rf<2><25> , \rf<2><24> ,
         \rf<2><23> , \rf<2><22> , \rf<2><21> , \rf<2><20> , \rf<2><19> ,
         \rf<2><18> , \rf<2><17> , \rf<2><16> , \rf<2><15> , \rf<2><14> ,
         \rf<2><13> , \rf<2><12> , \rf<2><11> , \rf<2><10> , \rf<2><9> ,
         \rf<2><8> , \rf<2><7> , \rf<2><6> , \rf<2><5> , \rf<2><4> ,
         \rf<2><3> , \rf<2><2> , \rf<2><1> , \rf<2><0> , \rf<1><31> ,
         \rf<1><30> , \rf<1><29> , \rf<1><28> , \rf<1><27> , \rf<1><26> ,
         \rf<1><25> , \rf<1><24> , \rf<1><23> , \rf<1><22> , \rf<1><21> ,
         \rf<1><20> , \rf<1><19> , \rf<1><18> , \rf<1><17> , \rf<1><16> ,
         \rf<1><15> , \rf<1><14> , \rf<1><13> , \rf<1><12> , \rf<1><11> ,
         \rf<1><10> , \rf<1><9> , \rf<1><8> , \rf<1><7> , \rf<1><6> ,
         \rf<1><5> , \rf<1><4> , \rf<1><3> , \rf<1><2> , \rf<1><1> ,
         \rf<1><0> , \rf<0><31> , \rf<0><30> , \rf<0><29> , \rf<0><28> ,
         \rf<0><27> , \rf<0><26> , \rf<0><25> , \rf<0><24> , \rf<0><23> ,
         \rf<0><22> , \rf<0><21> , \rf<0><20> , \rf<0><19> , \rf<0><18> ,
         \rf<0><17> , \rf<0><16> , \rf<0><15> , \rf<0><14> , \rf<0><13> ,
         \rf<0><12> , \rf<0><11> , \rf<0><10> , \rf<0><9> , \rf<0><8> ,
         \rf<0><7> , \rf<0><6> , \rf<0><5> , \rf<0><4> , \rf<0><3> ,
         \rf<0><2> , \rf<0><1> , \rf<0><0> , N503, N504, N505, N506, N507,
         N508, N509, N510, N511, N512, N513, N514, N515, N516, N517, N518,
         N519, N520, N521, N522, N523, N524, N525, N526, N527, N528, N529,
         N530, N531, N532, N533, N534, N536, N537, N538, N539, N540, N541,
         N542, N543, N544, N545, N546, N547, N548, N549, N550, N551, N552,
         N553, N554, N555, N556, N557, N558, N559, N560, N561, N562, N563,
         N564, N565, N566, N567, n534, n535, n537, n539, n541, n543, n548,
         n553, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28,
         n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42,
         n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56,
         n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84,
         n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98,
         n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
         n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763,
         n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774,
         n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785,
         n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796,
         n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807,
         n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818,
         n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829,
         n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840,
         n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851,
         n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862,
         n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873,
         n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884,
         n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895,
         n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906,
         n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917,
         n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928,
         n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939,
         n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950,
         n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961,
         n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972,
         n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983,
         n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994,
         n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
         n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
         n1045, n1046, n1047, n1048, n1049, n1050;
  assign N12 = \ra1<0> ;
  assign N13 = \ra1<1> ;
  assign N14 = \ra1<2> ;
  assign N15 = \ra1<3> ;
  assign N16 = \ra2<0> ;
  assign N17 = \ra2<1> ;
  assign N18 = \ra2<2> ;
  assign N19 = \ra2<3> ;

  EDFFXL \rf_reg<14><31>  ( .D(n5), .E(n977), .CK(clk), .Q(\rf<14><31> ) );
  EDFFXL \rf_reg<14><30>  ( .D(n975), .E(n977), .CK(clk), .Q(\rf<14><30> ) );
  EDFFXL \rf_reg<14><29>  ( .D(n2), .E(n977), .CK(clk), .Q(\rf<14><29> ) );
  EDFFXL \rf_reg<14><28>  ( .D(n1), .E(n977), .CK(clk), .Q(\rf<14><28> ) );
  EDFFXL \rf_reg<14><27>  ( .D(n972), .E(n977), .CK(clk), .Q(\rf<14><27> ) );
  EDFFXL \rf_reg<14><26>  ( .D(n971), .E(n977), .CK(clk), .Q(\rf<14><26> ) );
  EDFFXL \rf_reg<14><25>  ( .D(n970), .E(n977), .CK(clk), .Q(\rf<14><25> ) );
  EDFFXL \rf_reg<14><24>  ( .D(n969), .E(n19), .CK(clk), .Q(\rf<14><24> ) );
  EDFFXL \rf_reg<14><23>  ( .D(\wd3<23> ), .E(n19), .CK(clk), .Q(\rf<14><23> )
         );
  EDFFXL \rf_reg<14><22>  ( .D(n968), .E(n19), .CK(clk), .Q(\rf<14><22> ) );
  EDFFXL \rf_reg<14><21>  ( .D(n967), .E(n19), .CK(clk), .Q(\rf<14><21> ) );
  EDFFXL \rf_reg<14><20>  ( .D(n966), .E(n977), .CK(clk), .Q(\rf<14><20> ) );
  EDFFXL \rf_reg<14><19>  ( .D(n965), .E(n977), .CK(clk), .Q(\rf<14><19> ) );
  EDFFXL \rf_reg<14><18>  ( .D(n964), .E(n977), .CK(clk), .Q(\rf<14><18> ) );
  EDFFXL \rf_reg<14><17>  ( .D(n963), .E(n977), .CK(clk), .Q(\rf<14><17> ) );
  EDFFXL \rf_reg<14><16>  ( .D(n962), .E(n977), .CK(clk), .Q(\rf<14><16> ) );
  EDFFXL \rf_reg<14><15>  ( .D(\wd3<15> ), .E(n977), .CK(clk), .Q(\rf<14><15> ) );
  EDFFXL \rf_reg<14><14>  ( .D(\wd3<14> ), .E(n977), .CK(clk), .Q(\rf<14><14> ) );
  EDFFXL \rf_reg<14><13>  ( .D(\wd3<13> ), .E(n977), .CK(clk), .Q(\rf<14><13> ) );
  EDFFXL \rf_reg<14><12>  ( .D(\wd3<12> ), .E(n977), .CK(clk), .Q(\rf<14><12> ) );
  EDFFXL \rf_reg<14><11>  ( .D(n961), .E(n977), .CK(clk), .Q(\rf<14><11> ) );
  EDFFXL \rf_reg<14><10>  ( .D(n960), .E(n977), .CK(clk), .Q(\rf<14><10> ) );
  EDFFXL \rf_reg<14><9>  ( .D(n959), .E(n977), .CK(clk), .Q(\rf<14><9> ) );
  EDFFXL \rf_reg<14><8>  ( .D(n958), .E(n977), .CK(clk), .Q(\rf<14><8> ) );
  EDFFXL \rf_reg<14><7>  ( .D(n957), .E(n19), .CK(clk), .Q(\rf<14><7> ) );
  EDFFXL \rf_reg<14><6>  ( .D(n956), .E(n19), .CK(clk), .Q(\rf<14><6> ) );
  EDFFXL \rf_reg<14><5>  ( .D(n955), .E(n19), .CK(clk), .Q(\rf<14><5> ) );
  EDFFXL \rf_reg<14><4>  ( .D(n954), .E(n19), .CK(clk), .Q(\rf<14><4> ) );
  EDFFXL \rf_reg<14><3>  ( .D(n953), .E(n19), .CK(clk), .Q(\rf<14><3> ) );
  EDFFXL \rf_reg<14><2>  ( .D(n952), .E(n19), .CK(clk), .Q(\rf<14><2> ) );
  EDFFXL \rf_reg<14><1>  ( .D(n951), .E(n19), .CK(clk), .Q(\rf<14><1> ) );
  EDFFXL \rf_reg<14><0>  ( .D(n950), .E(n19), .CK(clk), .Q(\rf<14><0> ) );
  EDFFXL \rf_reg<13><31>  ( .D(n5), .E(n8), .CK(clk), .Q(\rf<13><31> ) );
  EDFFXL \rf_reg<13><30>  ( .D(n975), .E(n8), .CK(clk), .Q(\rf<13><30> ) );
  EDFFXL \rf_reg<13><29>  ( .D(n2), .E(n8), .CK(clk), .Q(\rf<13><29> ) );
  EDFFXL \rf_reg<13><28>  ( .D(n1), .E(n8), .CK(clk), .Q(\rf<13><28> ) );
  EDFFXL \rf_reg<13><27>  ( .D(n972), .E(n8), .CK(clk), .Q(\rf<13><27> ) );
  EDFFXL \rf_reg<13><26>  ( .D(n971), .E(n8), .CK(clk), .Q(\rf<13><26> ) );
  EDFFXL \rf_reg<13><25>  ( .D(n970), .E(n8), .CK(clk), .Q(\rf<13><25> ) );
  EDFFXL \rf_reg<13><24>  ( .D(n969), .E(n979), .CK(clk), .Q(\rf<13><24> ) );
  EDFFXL \rf_reg<13><23>  ( .D(\wd3<23> ), .E(n8), .CK(clk), .Q(\rf<13><23> )
         );
  EDFFXL \rf_reg<13><22>  ( .D(n968), .E(n8), .CK(clk), .Q(\rf<13><22> ) );
  EDFFXL \rf_reg<13><21>  ( .D(n967), .E(n8), .CK(clk), .Q(\rf<13><21> ) );
  EDFFXL \rf_reg<13><20>  ( .D(n966), .E(n979), .CK(clk), .Q(\rf<13><20> ) );
  EDFFXL \rf_reg<13><19>  ( .D(n965), .E(n979), .CK(clk), .Q(\rf<13><19> ) );
  EDFFXL \rf_reg<13><18>  ( .D(n964), .E(n979), .CK(clk), .Q(\rf<13><18> ) );
  EDFFXL \rf_reg<13><17>  ( .D(n963), .E(n979), .CK(clk), .Q(\rf<13><17> ) );
  EDFFXL \rf_reg<13><16>  ( .D(n962), .E(n979), .CK(clk), .Q(\rf<13><16> ) );
  EDFFXL \rf_reg<13><15>  ( .D(\wd3<15> ), .E(n979), .CK(clk), .Q(\rf<13><15> ) );
  EDFFXL \rf_reg<13><14>  ( .D(\wd3<14> ), .E(n979), .CK(clk), .Q(\rf<13><14> ) );
  EDFFXL \rf_reg<13><13>  ( .D(\wd3<13> ), .E(n979), .CK(clk), .Q(\rf<13><13> ) );
  EDFFXL \rf_reg<13><12>  ( .D(\wd3<12> ), .E(n979), .CK(clk), .Q(\rf<13><12> ) );
  EDFFXL \rf_reg<13><11>  ( .D(n961), .E(n979), .CK(clk), .Q(\rf<13><11> ) );
  EDFFXL \rf_reg<13><10>  ( .D(n960), .E(n979), .CK(clk), .Q(\rf<13><10> ) );
  EDFFXL \rf_reg<13><9>  ( .D(n959), .E(n979), .CK(clk), .Q(\rf<13><9> ) );
  EDFFXL \rf_reg<13><8>  ( .D(n958), .E(n979), .CK(clk), .Q(\rf<13><8> ) );
  EDFFXL \rf_reg<13><7>  ( .D(n957), .E(n979), .CK(clk), .Q(\rf<13><7> ) );
  EDFFXL \rf_reg<13><6>  ( .D(n956), .E(n979), .CK(clk), .Q(\rf<13><6> ) );
  EDFFXL \rf_reg<13><5>  ( .D(n955), .E(n979), .CK(clk), .Q(\rf<13><5> ) );
  EDFFXL \rf_reg<13><4>  ( .D(n954), .E(n979), .CK(clk), .Q(\rf<13><4> ) );
  EDFFXL \rf_reg<13><3>  ( .D(n953), .E(n979), .CK(clk), .Q(\rf<13><3> ) );
  EDFFXL \rf_reg<13><2>  ( .D(n952), .E(n979), .CK(clk), .Q(\rf<13><2> ) );
  EDFFXL \rf_reg<13><1>  ( .D(n951), .E(n8), .CK(clk), .Q(\rf<13><1> ) );
  EDFFXL \rf_reg<13><0>  ( .D(n950), .E(n8), .CK(clk), .Q(\rf<13><0> ) );
  EDFFXL \rf_reg<9><31>  ( .D(n5), .E(n7), .CK(clk), .Q(\rf<9><31> ) );
  EDFFXL \rf_reg<9><30>  ( .D(n975), .E(n7), .CK(clk), .Q(\rf<9><30> ) );
  EDFFXL \rf_reg<9><29>  ( .D(n2), .E(n7), .CK(clk), .Q(\rf<9><29> ) );
  EDFFXL \rf_reg<9><28>  ( .D(n1), .E(n7), .CK(clk), .Q(\rf<9><28> ) );
  EDFFXL \rf_reg<9><27>  ( .D(n972), .E(n7), .CK(clk), .Q(\rf<9><27> ) );
  EDFFXL \rf_reg<9><26>  ( .D(n971), .E(n7), .CK(clk), .Q(\rf<9><26> ) );
  EDFFXL \rf_reg<9><25>  ( .D(n970), .E(n7), .CK(clk), .Q(\rf<9><25> ) );
  EDFFXL \rf_reg<9><24>  ( .D(n969), .E(n987), .CK(clk), .Q(\rf<9><24> ) );
  EDFFXL \rf_reg<9><23>  ( .D(\wd3<23> ), .E(n7), .CK(clk), .Q(\rf<9><23> ) );
  EDFFXL \rf_reg<9><22>  ( .D(n968), .E(n7), .CK(clk), .Q(\rf<9><22> ) );
  EDFFXL \rf_reg<9><21>  ( .D(n967), .E(n7), .CK(clk), .Q(\rf<9><21> ) );
  EDFFXL \rf_reg<9><20>  ( .D(n966), .E(n987), .CK(clk), .Q(\rf<9><20> ) );
  EDFFXL \rf_reg<9><19>  ( .D(n965), .E(n987), .CK(clk), .Q(\rf<9><19> ) );
  EDFFXL \rf_reg<9><18>  ( .D(n964), .E(n987), .CK(clk), .Q(\rf<9><18> ) );
  EDFFXL \rf_reg<9><17>  ( .D(n963), .E(n987), .CK(clk), .Q(\rf<9><17> ) );
  EDFFXL \rf_reg<9><16>  ( .D(n962), .E(n987), .CK(clk), .Q(\rf<9><16> ) );
  EDFFXL \rf_reg<9><15>  ( .D(\wd3<15> ), .E(n987), .CK(clk), .Q(\rf<9><15> )
         );
  EDFFXL \rf_reg<9><14>  ( .D(\wd3<14> ), .E(n987), .CK(clk), .Q(\rf<9><14> )
         );
  EDFFXL \rf_reg<9><13>  ( .D(\wd3<13> ), .E(n987), .CK(clk), .Q(\rf<9><13> )
         );
  EDFFXL \rf_reg<9><12>  ( .D(\wd3<12> ), .E(n987), .CK(clk), .Q(\rf<9><12> )
         );
  EDFFXL \rf_reg<9><11>  ( .D(n961), .E(n987), .CK(clk), .Q(\rf<9><11> ) );
  EDFFXL \rf_reg<9><10>  ( .D(n960), .E(n987), .CK(clk), .Q(\rf<9><10> ) );
  EDFFXL \rf_reg<9><9>  ( .D(n959), .E(n987), .CK(clk), .Q(\rf<9><9> ) );
  EDFFXL \rf_reg<9><8>  ( .D(n958), .E(n987), .CK(clk), .Q(\rf<9><8> ) );
  EDFFXL \rf_reg<9><7>  ( .D(n957), .E(n987), .CK(clk), .Q(\rf<9><7> ) );
  EDFFXL \rf_reg<9><6>  ( .D(n956), .E(n987), .CK(clk), .Q(\rf<9><6> ) );
  EDFFXL \rf_reg<9><5>  ( .D(n955), .E(n987), .CK(clk), .Q(\rf<9><5> ) );
  EDFFXL \rf_reg<9><4>  ( .D(n954), .E(n987), .CK(clk), .Q(\rf<9><4> ) );
  EDFFXL \rf_reg<9><3>  ( .D(n953), .E(n987), .CK(clk), .Q(\rf<9><3> ) );
  EDFFXL \rf_reg<9><2>  ( .D(n952), .E(n987), .CK(clk), .Q(\rf<9><2> ) );
  EDFFXL \rf_reg<9><1>  ( .D(n951), .E(n7), .CK(clk), .Q(\rf<9><1> ) );
  EDFFXL \rf_reg<9><0>  ( .D(n950), .E(n7), .CK(clk), .Q(\rf<9><0> ) );
  EDFFXL \rf_reg<5><31>  ( .D(n5), .E(n995), .CK(clk), .Q(\rf<5><31> ) );
  EDFFXL \rf_reg<5><30>  ( .D(n975), .E(n995), .CK(clk), .Q(\rf<5><30> ) );
  EDFFXL \rf_reg<5><29>  ( .D(n2), .E(n995), .CK(clk), .Q(\rf<5><29> ) );
  EDFFXL \rf_reg<5><28>  ( .D(n1), .E(n995), .CK(clk), .Q(\rf<5><28> ) );
  EDFFXL \rf_reg<5><27>  ( .D(n972), .E(n995), .CK(clk), .Q(\rf<5><27> ) );
  EDFFXL \rf_reg<5><26>  ( .D(n971), .E(n995), .CK(clk), .Q(\rf<5><26> ) );
  EDFFXL \rf_reg<5><25>  ( .D(n970), .E(n995), .CK(clk), .Q(\rf<5><25> ) );
  EDFFXL \rf_reg<5><24>  ( .D(n969), .E(n6), .CK(clk), .Q(\rf<5><24> ) );
  EDFFXL \rf_reg<5><23>  ( .D(\wd3<23> ), .E(n6), .CK(clk), .Q(\rf<5><23> ) );
  EDFFXL \rf_reg<5><22>  ( .D(n968), .E(n6), .CK(clk), .Q(\rf<5><22> ) );
  EDFFXL \rf_reg<5><21>  ( .D(n967), .E(n6), .CK(clk), .Q(\rf<5><21> ) );
  EDFFXL \rf_reg<5><20>  ( .D(n966), .E(n995), .CK(clk), .Q(\rf<5><20> ) );
  EDFFXL \rf_reg<5><19>  ( .D(n965), .E(n995), .CK(clk), .Q(\rf<5><19> ) );
  EDFFXL \rf_reg<5><18>  ( .D(n964), .E(n995), .CK(clk), .Q(\rf<5><18> ) );
  EDFFXL \rf_reg<5><17>  ( .D(n963), .E(n995), .CK(clk), .Q(\rf<5><17> ) );
  EDFFXL \rf_reg<5><16>  ( .D(n962), .E(n995), .CK(clk), .Q(\rf<5><16> ) );
  EDFFXL \rf_reg<5><15>  ( .D(\wd3<15> ), .E(n995), .CK(clk), .Q(\rf<5><15> )
         );
  EDFFXL \rf_reg<5><14>  ( .D(\wd3<14> ), .E(n995), .CK(clk), .Q(\rf<5><14> )
         );
  EDFFXL \rf_reg<5><13>  ( .D(\wd3<13> ), .E(n995), .CK(clk), .Q(\rf<5><13> )
         );
  EDFFXL \rf_reg<5><12>  ( .D(\wd3<12> ), .E(n995), .CK(clk), .Q(\rf<5><12> )
         );
  EDFFXL \rf_reg<5><11>  ( .D(n961), .E(n995), .CK(clk), .Q(\rf<5><11> ) );
  EDFFXL \rf_reg<5><10>  ( .D(n960), .E(n995), .CK(clk), .Q(\rf<5><10> ) );
  EDFFXL \rf_reg<5><9>  ( .D(n959), .E(n995), .CK(clk), .Q(\rf<5><9> ) );
  EDFFXL \rf_reg<5><8>  ( .D(n958), .E(n995), .CK(clk), .Q(\rf<5><8> ) );
  EDFFXL \rf_reg<5><7>  ( .D(n957), .E(n6), .CK(clk), .Q(\rf<5><7> ) );
  EDFFXL \rf_reg<5><6>  ( .D(n956), .E(n6), .CK(clk), .Q(\rf<5><6> ) );
  EDFFXL \rf_reg<5><5>  ( .D(n955), .E(n6), .CK(clk), .Q(\rf<5><5> ) );
  EDFFXL \rf_reg<5><4>  ( .D(n954), .E(n6), .CK(clk), .Q(\rf<5><4> ) );
  EDFFXL \rf_reg<5><3>  ( .D(n953), .E(n6), .CK(clk), .Q(\rf<5><3> ) );
  EDFFXL \rf_reg<5><2>  ( .D(n952), .E(n6), .CK(clk), .Q(\rf<5><2> ) );
  EDFFXL \rf_reg<5><1>  ( .D(n951), .E(n6), .CK(clk), .Q(\rf<5><1> ) );
  EDFFXL \rf_reg<5><0>  ( .D(n950), .E(n6), .CK(clk), .Q(\rf<5><0> ) );
  EDFFXL \rf_reg<1><31>  ( .D(n5), .E(n1003), .CK(clk), .Q(\rf<1><31> ) );
  EDFFXL \rf_reg<1><30>  ( .D(n975), .E(n1003), .CK(clk), .Q(\rf<1><30> ) );
  EDFFXL \rf_reg<1><29>  ( .D(n2), .E(n1003), .CK(clk), .Q(\rf<1><29> ) );
  EDFFXL \rf_reg<1><28>  ( .D(n1), .E(n1003), .CK(clk), .Q(\rf<1><28> ) );
  EDFFXL \rf_reg<1><27>  ( .D(n972), .E(n1003), .CK(clk), .Q(\rf<1><27> ) );
  EDFFXL \rf_reg<1><26>  ( .D(n971), .E(n1003), .CK(clk), .Q(\rf<1><26> ) );
  EDFFXL \rf_reg<1><25>  ( .D(n970), .E(n1003), .CK(clk), .Q(\rf<1><25> ) );
  EDFFXL \rf_reg<1><24>  ( .D(n969), .E(n10), .CK(clk), .Q(\rf<1><24> ) );
  EDFFXL \rf_reg<1><23>  ( .D(\wd3<23> ), .E(n10), .CK(clk), .Q(\rf<1><23> )
         );
  EDFFXL \rf_reg<1><22>  ( .D(n968), .E(n10), .CK(clk), .Q(\rf<1><22> ) );
  EDFFXL \rf_reg<1><21>  ( .D(n967), .E(n10), .CK(clk), .Q(\rf<1><21> ) );
  EDFFXL \rf_reg<1><20>  ( .D(n966), .E(n1003), .CK(clk), .Q(\rf<1><20> ) );
  EDFFXL \rf_reg<1><19>  ( .D(n965), .E(n1003), .CK(clk), .Q(\rf<1><19> ) );
  EDFFXL \rf_reg<1><18>  ( .D(n964), .E(n1003), .CK(clk), .Q(\rf<1><18> ) );
  EDFFXL \rf_reg<1><17>  ( .D(n963), .E(n1003), .CK(clk), .Q(\rf<1><17> ) );
  EDFFXL \rf_reg<1><16>  ( .D(n962), .E(n1003), .CK(clk), .Q(\rf<1><16> ) );
  EDFFXL \rf_reg<1><15>  ( .D(\wd3<15> ), .E(n1003), .CK(clk), .Q(\rf<1><15> )
         );
  EDFFXL \rf_reg<1><14>  ( .D(\wd3<14> ), .E(n1003), .CK(clk), .Q(\rf<1><14> )
         );
  EDFFXL \rf_reg<1><13>  ( .D(\wd3<13> ), .E(n1003), .CK(clk), .Q(\rf<1><13> )
         );
  EDFFXL \rf_reg<1><12>  ( .D(\wd3<12> ), .E(n1003), .CK(clk), .Q(\rf<1><12> )
         );
  EDFFXL \rf_reg<1><11>  ( .D(n961), .E(n1003), .CK(clk), .Q(\rf<1><11> ) );
  EDFFXL \rf_reg<1><10>  ( .D(n960), .E(n1003), .CK(clk), .Q(\rf<1><10> ) );
  EDFFXL \rf_reg<1><9>  ( .D(n959), .E(n1003), .CK(clk), .Q(\rf<1><9> ) );
  EDFFXL \rf_reg<1><8>  ( .D(n958), .E(n1003), .CK(clk), .Q(\rf<1><8> ) );
  EDFFXL \rf_reg<1><7>  ( .D(n957), .E(n10), .CK(clk), .Q(\rf<1><7> ) );
  EDFFXL \rf_reg<1><6>  ( .D(n956), .E(n10), .CK(clk), .Q(\rf<1><6> ) );
  EDFFXL \rf_reg<1><5>  ( .D(n955), .E(n10), .CK(clk), .Q(\rf<1><5> ) );
  EDFFXL \rf_reg<1><4>  ( .D(n954), .E(n10), .CK(clk), .Q(\rf<1><4> ) );
  EDFFXL \rf_reg<1><3>  ( .D(n953), .E(n10), .CK(clk), .Q(\rf<1><3> ) );
  EDFFXL \rf_reg<1><2>  ( .D(n952), .E(n10), .CK(clk), .Q(\rf<1><2> ) );
  EDFFXL \rf_reg<1><1>  ( .D(n951), .E(n10), .CK(clk), .Q(\rf<1><1> ) );
  EDFFXL \rf_reg<1><0>  ( .D(n950), .E(n10), .CK(clk), .Q(\rf<1><0> ) );
  EDFFXL \rf_reg<11><31>  ( .D(n5), .E(n983), .CK(clk), .Q(\rf<11><31> ) );
  EDFFXL \rf_reg<11><30>  ( .D(n975), .E(n983), .CK(clk), .Q(\rf<11><30> ) );
  EDFFXL \rf_reg<11><29>  ( .D(n2), .E(n983), .CK(clk), .Q(\rf<11><29> ) );
  EDFFXL \rf_reg<11><28>  ( .D(n1), .E(n983), .CK(clk), .Q(\rf<11><28> ) );
  EDFFXL \rf_reg<11><27>  ( .D(n972), .E(n983), .CK(clk), .Q(\rf<11><27> ) );
  EDFFXL \rf_reg<11><26>  ( .D(n971), .E(n983), .CK(clk), .Q(\rf<11><26> ) );
  EDFFXL \rf_reg<11><25>  ( .D(n970), .E(n983), .CK(clk), .Q(\rf<11><25> ) );
  EDFFXL \rf_reg<11><24>  ( .D(n969), .E(n20), .CK(clk), .Q(\rf<11><24> ) );
  EDFFXL \rf_reg<11><23>  ( .D(\wd3<23> ), .E(n20), .CK(clk), .Q(\rf<11><23> )
         );
  EDFFXL \rf_reg<11><22>  ( .D(n968), .E(n20), .CK(clk), .Q(\rf<11><22> ) );
  EDFFXL \rf_reg<11><21>  ( .D(n967), .E(n20), .CK(clk), .Q(\rf<11><21> ) );
  EDFFXL \rf_reg<11><20>  ( .D(n966), .E(n983), .CK(clk), .Q(\rf<11><20> ) );
  EDFFXL \rf_reg<11><19>  ( .D(n965), .E(n983), .CK(clk), .Q(\rf<11><19> ) );
  EDFFXL \rf_reg<11><18>  ( .D(n964), .E(n983), .CK(clk), .Q(\rf<11><18> ) );
  EDFFXL \rf_reg<11><17>  ( .D(n963), .E(n983), .CK(clk), .Q(\rf<11><17> ) );
  EDFFXL \rf_reg<11><16>  ( .D(n962), .E(n983), .CK(clk), .Q(\rf<11><16> ) );
  EDFFXL \rf_reg<11><15>  ( .D(\wd3<15> ), .E(n983), .CK(clk), .Q(\rf<11><15> ) );
  EDFFXL \rf_reg<11><14>  ( .D(\wd3<14> ), .E(n983), .CK(clk), .Q(\rf<11><14> ) );
  EDFFXL \rf_reg<11><13>  ( .D(\wd3<13> ), .E(n983), .CK(clk), .Q(\rf<11><13> ) );
  EDFFXL \rf_reg<11><12>  ( .D(\wd3<12> ), .E(n983), .CK(clk), .Q(\rf<11><12> ) );
  EDFFXL \rf_reg<11><11>  ( .D(n961), .E(n983), .CK(clk), .Q(\rf<11><11> ) );
  EDFFXL \rf_reg<11><10>  ( .D(n960), .E(n983), .CK(clk), .Q(\rf<11><10> ) );
  EDFFXL \rf_reg<11><9>  ( .D(n959), .E(n983), .CK(clk), .Q(\rf<11><9> ) );
  EDFFXL \rf_reg<11><8>  ( .D(n958), .E(n983), .CK(clk), .Q(\rf<11><8> ) );
  EDFFXL \rf_reg<11><7>  ( .D(n957), .E(n20), .CK(clk), .Q(\rf<11><7> ) );
  EDFFXL \rf_reg<11><6>  ( .D(n956), .E(n20), .CK(clk), .Q(\rf<11><6> ) );
  EDFFXL \rf_reg<11><5>  ( .D(n955), .E(n20), .CK(clk), .Q(\rf<11><5> ) );
  EDFFXL \rf_reg<11><4>  ( .D(n954), .E(n20), .CK(clk), .Q(\rf<11><4> ) );
  EDFFXL \rf_reg<11><3>  ( .D(n953), .E(n20), .CK(clk), .Q(\rf<11><3> ) );
  EDFFXL \rf_reg<11><2>  ( .D(n952), .E(n20), .CK(clk), .Q(\rf<11><2> ) );
  EDFFXL \rf_reg<11><1>  ( .D(n951), .E(n20), .CK(clk), .Q(\rf<11><1> ) );
  EDFFXL \rf_reg<11><0>  ( .D(n950), .E(n20), .CK(clk), .Q(\rf<11><0> ) );
  EDFFXL \rf_reg<7><31>  ( .D(n5), .E(n991), .CK(clk), .Q(\rf<7><31> ) );
  EDFFXL \rf_reg<7><30>  ( .D(n975), .E(n991), .CK(clk), .Q(\rf<7><30> ) );
  EDFFXL \rf_reg<7><29>  ( .D(n2), .E(n991), .CK(clk), .Q(\rf<7><29> ) );
  EDFFXL \rf_reg<7><28>  ( .D(n1), .E(n991), .CK(clk), .Q(\rf<7><28> ) );
  EDFFXL \rf_reg<7><27>  ( .D(n972), .E(n991), .CK(clk), .Q(\rf<7><27> ) );
  EDFFXL \rf_reg<7><26>  ( .D(n971), .E(n991), .CK(clk), .Q(\rf<7><26> ) );
  EDFFXL \rf_reg<7><25>  ( .D(n970), .E(n991), .CK(clk), .Q(\rf<7><25> ) );
  EDFFXL \rf_reg<7><24>  ( .D(n969), .E(n17), .CK(clk), .Q(\rf<7><24> ) );
  EDFFXL \rf_reg<7><23>  ( .D(\wd3<23> ), .E(n17), .CK(clk), .Q(\rf<7><23> )
         );
  EDFFXL \rf_reg<7><22>  ( .D(n968), .E(n17), .CK(clk), .Q(\rf<7><22> ) );
  EDFFXL \rf_reg<7><21>  ( .D(n967), .E(n17), .CK(clk), .Q(\rf<7><21> ) );
  EDFFXL \rf_reg<7><20>  ( .D(n966), .E(n991), .CK(clk), .Q(\rf<7><20> ) );
  EDFFXL \rf_reg<7><19>  ( .D(n965), .E(n991), .CK(clk), .Q(\rf<7><19> ) );
  EDFFXL \rf_reg<7><18>  ( .D(n964), .E(n991), .CK(clk), .Q(\rf<7><18> ) );
  EDFFXL \rf_reg<7><17>  ( .D(n963), .E(n991), .CK(clk), .Q(\rf<7><17> ) );
  EDFFXL \rf_reg<7><16>  ( .D(n962), .E(n991), .CK(clk), .Q(\rf<7><16> ) );
  EDFFXL \rf_reg<7><15>  ( .D(\wd3<15> ), .E(n991), .CK(clk), .Q(\rf<7><15> )
         );
  EDFFXL \rf_reg<7><14>  ( .D(\wd3<14> ), .E(n991), .CK(clk), .Q(\rf<7><14> )
         );
  EDFFXL \rf_reg<7><13>  ( .D(\wd3<13> ), .E(n991), .CK(clk), .Q(\rf<7><13> )
         );
  EDFFXL \rf_reg<7><12>  ( .D(\wd3<12> ), .E(n991), .CK(clk), .Q(\rf<7><12> )
         );
  EDFFXL \rf_reg<7><11>  ( .D(n961), .E(n991), .CK(clk), .Q(\rf<7><11> ) );
  EDFFXL \rf_reg<7><10>  ( .D(n960), .E(n991), .CK(clk), .Q(\rf<7><10> ) );
  EDFFXL \rf_reg<7><9>  ( .D(n959), .E(n991), .CK(clk), .Q(\rf<7><9> ) );
  EDFFXL \rf_reg<7><8>  ( .D(n958), .E(n991), .CK(clk), .Q(\rf<7><8> ) );
  EDFFXL \rf_reg<7><7>  ( .D(n957), .E(n17), .CK(clk), .Q(\rf<7><7> ) );
  EDFFXL \rf_reg<7><6>  ( .D(n956), .E(n17), .CK(clk), .Q(\rf<7><6> ) );
  EDFFXL \rf_reg<7><5>  ( .D(n955), .E(n17), .CK(clk), .Q(\rf<7><5> ) );
  EDFFXL \rf_reg<7><4>  ( .D(n954), .E(n17), .CK(clk), .Q(\rf<7><4> ) );
  EDFFXL \rf_reg<7><3>  ( .D(n953), .E(n17), .CK(clk), .Q(\rf<7><3> ) );
  EDFFXL \rf_reg<7><2>  ( .D(n952), .E(n17), .CK(clk), .Q(\rf<7><2> ) );
  EDFFXL \rf_reg<7><1>  ( .D(n951), .E(n17), .CK(clk), .Q(\rf<7><1> ) );
  EDFFXL \rf_reg<7><0>  ( .D(n950), .E(n17), .CK(clk), .Q(\rf<7><0> ) );
  EDFFXL \rf_reg<3><31>  ( .D(n5), .E(n999), .CK(clk), .Q(\rf<3><31> ) );
  EDFFXL \rf_reg<3><30>  ( .D(n975), .E(n999), .CK(clk), .Q(\rf<3><30> ) );
  EDFFXL \rf_reg<3><29>  ( .D(n2), .E(n999), .CK(clk), .Q(\rf<3><29> ) );
  EDFFXL \rf_reg<3><28>  ( .D(n1), .E(n999), .CK(clk), .Q(\rf<3><28> ) );
  EDFFXL \rf_reg<3><27>  ( .D(n972), .E(n999), .CK(clk), .Q(\rf<3><27> ) );
  EDFFXL \rf_reg<3><26>  ( .D(n971), .E(n999), .CK(clk), .Q(\rf<3><26> ) );
  EDFFXL \rf_reg<3><25>  ( .D(n970), .E(n999), .CK(clk), .Q(\rf<3><25> ) );
  EDFFXL \rf_reg<3><24>  ( .D(n969), .E(n12), .CK(clk), .Q(\rf<3><24> ) );
  EDFFXL \rf_reg<3><23>  ( .D(\wd3<23> ), .E(n12), .CK(clk), .Q(\rf<3><23> )
         );
  EDFFXL \rf_reg<3><22>  ( .D(n968), .E(n12), .CK(clk), .Q(\rf<3><22> ) );
  EDFFXL \rf_reg<3><21>  ( .D(n967), .E(n12), .CK(clk), .Q(\rf<3><21> ) );
  EDFFXL \rf_reg<3><20>  ( .D(n966), .E(n999), .CK(clk), .Q(\rf<3><20> ) );
  EDFFXL \rf_reg<3><19>  ( .D(n965), .E(n999), .CK(clk), .Q(\rf<3><19> ) );
  EDFFXL \rf_reg<3><18>  ( .D(n964), .E(n999), .CK(clk), .Q(\rf<3><18> ) );
  EDFFXL \rf_reg<3><17>  ( .D(n963), .E(n999), .CK(clk), .Q(\rf<3><17> ) );
  EDFFXL \rf_reg<3><16>  ( .D(n962), .E(n999), .CK(clk), .Q(\rf<3><16> ) );
  EDFFXL \rf_reg<3><15>  ( .D(\wd3<15> ), .E(n999), .CK(clk), .Q(\rf<3><15> )
         );
  EDFFXL \rf_reg<3><14>  ( .D(\wd3<14> ), .E(n999), .CK(clk), .Q(\rf<3><14> )
         );
  EDFFXL \rf_reg<3><13>  ( .D(\wd3<13> ), .E(n999), .CK(clk), .Q(\rf<3><13> )
         );
  EDFFXL \rf_reg<3><12>  ( .D(\wd3<12> ), .E(n999), .CK(clk), .Q(\rf<3><12> )
         );
  EDFFXL \rf_reg<3><11>  ( .D(n961), .E(n999), .CK(clk), .Q(\rf<3><11> ) );
  EDFFXL \rf_reg<3><10>  ( .D(n960), .E(n999), .CK(clk), .Q(\rf<3><10> ) );
  EDFFXL \rf_reg<3><9>  ( .D(n959), .E(n999), .CK(clk), .Q(\rf<3><9> ) );
  EDFFXL \rf_reg<3><8>  ( .D(n958), .E(n999), .CK(clk), .Q(\rf<3><8> ) );
  EDFFXL \rf_reg<3><7>  ( .D(n957), .E(n12), .CK(clk), .Q(\rf<3><7> ) );
  EDFFXL \rf_reg<3><6>  ( .D(n956), .E(n12), .CK(clk), .Q(\rf<3><6> ) );
  EDFFXL \rf_reg<3><5>  ( .D(n955), .E(n12), .CK(clk), .Q(\rf<3><5> ) );
  EDFFXL \rf_reg<3><4>  ( .D(n954), .E(n12), .CK(clk), .Q(\rf<3><4> ) );
  EDFFXL \rf_reg<3><3>  ( .D(n953), .E(n12), .CK(clk), .Q(\rf<3><3> ) );
  EDFFXL \rf_reg<3><2>  ( .D(n952), .E(n12), .CK(clk), .Q(\rf<3><2> ) );
  EDFFXL \rf_reg<3><1>  ( .D(n951), .E(n12), .CK(clk), .Q(\rf<3><1> ) );
  EDFFXL \rf_reg<3><0>  ( .D(n950), .E(n12), .CK(clk), .Q(\rf<3><0> ) );
  EDFFXL \rf_reg<8><31>  ( .D(n5), .E(n989), .CK(clk), .Q(\rf<8><31> ) );
  EDFFXL \rf_reg<8><30>  ( .D(n975), .E(n989), .CK(clk), .Q(\rf<8><30> ) );
  EDFFXL \rf_reg<8><29>  ( .D(n2), .E(n989), .CK(clk), .Q(\rf<8><29> ) );
  EDFFXL \rf_reg<8><28>  ( .D(n1), .E(n989), .CK(clk), .Q(\rf<8><28> ) );
  EDFFXL \rf_reg<8><27>  ( .D(n972), .E(n989), .CK(clk), .Q(\rf<8><27> ) );
  EDFFXL \rf_reg<8><26>  ( .D(n971), .E(n989), .CK(clk), .Q(\rf<8><26> ) );
  EDFFXL \rf_reg<8><25>  ( .D(n970), .E(n989), .CK(clk), .Q(\rf<8><25> ) );
  EDFFXL \rf_reg<8><24>  ( .D(n969), .E(n14), .CK(clk), .Q(\rf<8><24> ) );
  EDFFXL \rf_reg<8><23>  ( .D(\wd3<23> ), .E(n14), .CK(clk), .Q(\rf<8><23> )
         );
  EDFFXL \rf_reg<8><22>  ( .D(n968), .E(n14), .CK(clk), .Q(\rf<8><22> ) );
  EDFFXL \rf_reg<8><21>  ( .D(n967), .E(n14), .CK(clk), .Q(\rf<8><21> ) );
  EDFFXL \rf_reg<8><20>  ( .D(n966), .E(n989), .CK(clk), .Q(\rf<8><20> ) );
  EDFFXL \rf_reg<8><19>  ( .D(n965), .E(n989), .CK(clk), .Q(\rf<8><19> ) );
  EDFFXL \rf_reg<8><18>  ( .D(n964), .E(n989), .CK(clk), .Q(\rf<8><18> ) );
  EDFFXL \rf_reg<8><17>  ( .D(n963), .E(n989), .CK(clk), .Q(\rf<8><17> ) );
  EDFFXL \rf_reg<8><16>  ( .D(n962), .E(n989), .CK(clk), .Q(\rf<8><16> ) );
  EDFFXL \rf_reg<8><15>  ( .D(\wd3<15> ), .E(n989), .CK(clk), .Q(\rf<8><15> )
         );
  EDFFXL \rf_reg<8><14>  ( .D(\wd3<14> ), .E(n989), .CK(clk), .Q(\rf<8><14> )
         );
  EDFFXL \rf_reg<8><13>  ( .D(\wd3<13> ), .E(n989), .CK(clk), .Q(\rf<8><13> )
         );
  EDFFXL \rf_reg<8><12>  ( .D(\wd3<12> ), .E(n989), .CK(clk), .Q(\rf<8><12> )
         );
  EDFFXL \rf_reg<8><11>  ( .D(n961), .E(n989), .CK(clk), .Q(\rf<8><11> ) );
  EDFFXL \rf_reg<8><10>  ( .D(n960), .E(n989), .CK(clk), .Q(\rf<8><10> ) );
  EDFFXL \rf_reg<8><9>  ( .D(n959), .E(n989), .CK(clk), .Q(\rf<8><9> ) );
  EDFFXL \rf_reg<8><8>  ( .D(n958), .E(n989), .CK(clk), .Q(\rf<8><8> ) );
  EDFFXL \rf_reg<8><7>  ( .D(n957), .E(n14), .CK(clk), .Q(\rf<8><7> ) );
  EDFFXL \rf_reg<8><6>  ( .D(n956), .E(n14), .CK(clk), .Q(\rf<8><6> ) );
  EDFFXL \rf_reg<8><5>  ( .D(n955), .E(n14), .CK(clk), .Q(\rf<8><5> ) );
  EDFFXL \rf_reg<8><4>  ( .D(n954), .E(n14), .CK(clk), .Q(\rf<8><4> ) );
  EDFFXL \rf_reg<8><3>  ( .D(n953), .E(n14), .CK(clk), .Q(\rf<8><3> ) );
  EDFFXL \rf_reg<8><2>  ( .D(n952), .E(n14), .CK(clk), .Q(\rf<8><2> ) );
  EDFFXL \rf_reg<8><1>  ( .D(n951), .E(n14), .CK(clk), .Q(\rf<8><1> ) );
  EDFFXL \rf_reg<8><0>  ( .D(n950), .E(n14), .CK(clk), .Q(\rf<8><0> ) );
  EDFFXL \rf_reg<4><31>  ( .D(n5), .E(n997), .CK(clk), .Q(\rf<4><31> ) );
  EDFFXL \rf_reg<4><30>  ( .D(n975), .E(n997), .CK(clk), .Q(\rf<4><30> ) );
  EDFFXL \rf_reg<4><29>  ( .D(n2), .E(n997), .CK(clk), .Q(\rf<4><29> ) );
  EDFFXL \rf_reg<4><28>  ( .D(n1), .E(n997), .CK(clk), .Q(\rf<4><28> ) );
  EDFFXL \rf_reg<4><27>  ( .D(n972), .E(n997), .CK(clk), .Q(\rf<4><27> ) );
  EDFFXL \rf_reg<4><26>  ( .D(n971), .E(n997), .CK(clk), .Q(\rf<4><26> ) );
  EDFFXL \rf_reg<4><25>  ( .D(n970), .E(n997), .CK(clk), .Q(\rf<4><25> ) );
  EDFFXL \rf_reg<4><24>  ( .D(n969), .E(n13), .CK(clk), .Q(\rf<4><24> ) );
  EDFFXL \rf_reg<4><23>  ( .D(\wd3<23> ), .E(n13), .CK(clk), .Q(\rf<4><23> )
         );
  EDFFXL \rf_reg<4><22>  ( .D(n968), .E(n13), .CK(clk), .Q(\rf<4><22> ) );
  EDFFXL \rf_reg<4><21>  ( .D(n967), .E(n13), .CK(clk), .Q(\rf<4><21> ) );
  EDFFXL \rf_reg<4><20>  ( .D(n966), .E(n997), .CK(clk), .Q(\rf<4><20> ) );
  EDFFXL \rf_reg<4><19>  ( .D(n965), .E(n997), .CK(clk), .Q(\rf<4><19> ) );
  EDFFXL \rf_reg<4><18>  ( .D(n964), .E(n997), .CK(clk), .Q(\rf<4><18> ) );
  EDFFXL \rf_reg<4><17>  ( .D(n963), .E(n997), .CK(clk), .Q(\rf<4><17> ) );
  EDFFXL \rf_reg<4><16>  ( .D(n962), .E(n997), .CK(clk), .Q(\rf<4><16> ) );
  EDFFXL \rf_reg<4><15>  ( .D(\wd3<15> ), .E(n997), .CK(clk), .Q(\rf<4><15> )
         );
  EDFFXL \rf_reg<4><14>  ( .D(\wd3<14> ), .E(n997), .CK(clk), .Q(\rf<4><14> )
         );
  EDFFXL \rf_reg<4><13>  ( .D(\wd3<13> ), .E(n997), .CK(clk), .Q(\rf<4><13> )
         );
  EDFFXL \rf_reg<4><12>  ( .D(\wd3<12> ), .E(n997), .CK(clk), .Q(\rf<4><12> )
         );
  EDFFXL \rf_reg<4><11>  ( .D(n961), .E(n997), .CK(clk), .Q(\rf<4><11> ) );
  EDFFXL \rf_reg<4><10>  ( .D(n960), .E(n997), .CK(clk), .Q(\rf<4><10> ) );
  EDFFXL \rf_reg<4><9>  ( .D(n959), .E(n997), .CK(clk), .Q(\rf<4><9> ) );
  EDFFXL \rf_reg<4><8>  ( .D(n958), .E(n997), .CK(clk), .Q(\rf<4><8> ) );
  EDFFXL \rf_reg<4><7>  ( .D(n957), .E(n13), .CK(clk), .Q(\rf<4><7> ) );
  EDFFXL \rf_reg<4><6>  ( .D(n956), .E(n13), .CK(clk), .Q(\rf<4><6> ) );
  EDFFXL \rf_reg<4><5>  ( .D(n955), .E(n13), .CK(clk), .Q(\rf<4><5> ) );
  EDFFXL \rf_reg<4><4>  ( .D(n954), .E(n13), .CK(clk), .Q(\rf<4><4> ) );
  EDFFXL \rf_reg<4><3>  ( .D(n953), .E(n13), .CK(clk), .Q(\rf<4><3> ) );
  EDFFXL \rf_reg<4><2>  ( .D(n952), .E(n13), .CK(clk), .Q(\rf<4><2> ) );
  EDFFXL \rf_reg<4><1>  ( .D(n951), .E(n13), .CK(clk), .Q(\rf<4><1> ) );
  EDFFXL \rf_reg<4><0>  ( .D(n950), .E(n13), .CK(clk), .Q(\rf<4><0> ) );
  EDFFXL \rf_reg<0><31>  ( .D(n5), .E(n9), .CK(clk), .Q(\rf<0><31> ) );
  EDFFXL \rf_reg<0><30>  ( .D(n975), .E(n9), .CK(clk), .Q(\rf<0><30> ) );
  EDFFXL \rf_reg<0><29>  ( .D(n2), .E(n9), .CK(clk), .Q(\rf<0><29> ) );
  EDFFXL \rf_reg<0><28>  ( .D(n1), .E(n9), .CK(clk), .Q(\rf<0><28> ) );
  EDFFXL \rf_reg<0><27>  ( .D(n972), .E(n9), .CK(clk), .Q(\rf<0><27> ) );
  EDFFXL \rf_reg<0><26>  ( .D(n971), .E(n9), .CK(clk), .Q(\rf<0><26> ) );
  EDFFXL \rf_reg<0><25>  ( .D(n970), .E(n9), .CK(clk), .Q(\rf<0><25> ) );
  EDFFXL \rf_reg<0><24>  ( .D(n969), .E(n9), .CK(clk), .Q(\rf<0><24> ) );
  EDFFXL \rf_reg<0><23>  ( .D(\wd3<23> ), .E(n1005), .CK(clk), .Q(\rf<0><23> )
         );
  EDFFXL \rf_reg<0><22>  ( .D(n968), .E(n1005), .CK(clk), .Q(\rf<0><22> ) );
  EDFFXL \rf_reg<0><21>  ( .D(n967), .E(n1005), .CK(clk), .Q(\rf<0><21> ) );
  EDFFXL \rf_reg<0><20>  ( .D(n966), .E(n1005), .CK(clk), .Q(\rf<0><20> ) );
  EDFFXL \rf_reg<0><19>  ( .D(n965), .E(n1005), .CK(clk), .Q(\rf<0><19> ) );
  EDFFXL \rf_reg<0><18>  ( .D(n964), .E(n1005), .CK(clk), .Q(\rf<0><18> ) );
  EDFFXL \rf_reg<0><17>  ( .D(n963), .E(n1005), .CK(clk), .Q(\rf<0><17> ) );
  EDFFXL \rf_reg<0><16>  ( .D(n962), .E(n1005), .CK(clk), .Q(\rf<0><16> ) );
  EDFFXL \rf_reg<0><15>  ( .D(\wd3<15> ), .E(n1005), .CK(clk), .Q(\rf<0><15> )
         );
  EDFFXL \rf_reg<0><14>  ( .D(\wd3<14> ), .E(n1005), .CK(clk), .Q(\rf<0><14> )
         );
  EDFFXL \rf_reg<0><13>  ( .D(\wd3<13> ), .E(n1005), .CK(clk), .Q(\rf<0><13> )
         );
  EDFFXL \rf_reg<0><12>  ( .D(\wd3<12> ), .E(n9), .CK(clk), .Q(\rf<0><12> ) );
  EDFFXL \rf_reg<0><11>  ( .D(n961), .E(n9), .CK(clk), .Q(\rf<0><11> ) );
  EDFFXL \rf_reg<0><10>  ( .D(n960), .E(n9), .CK(clk), .Q(\rf<0><10> ) );
  EDFFXL \rf_reg<0><9>  ( .D(n959), .E(n9), .CK(clk), .Q(\rf<0><9> ) );
  EDFFXL \rf_reg<0><8>  ( .D(n958), .E(n1005), .CK(clk), .Q(\rf<0><8> ) );
  EDFFXL \rf_reg<0><7>  ( .D(n957), .E(n1005), .CK(clk), .Q(\rf<0><7> ) );
  EDFFXL \rf_reg<0><6>  ( .D(n956), .E(n1005), .CK(clk), .Q(\rf<0><6> ) );
  EDFFXL \rf_reg<0><5>  ( .D(n955), .E(n1005), .CK(clk), .Q(\rf<0><5> ) );
  EDFFXL \rf_reg<0><4>  ( .D(n954), .E(n1005), .CK(clk), .Q(\rf<0><4> ) );
  EDFFXL \rf_reg<0><3>  ( .D(n953), .E(n1005), .CK(clk), .Q(\rf<0><3> ) );
  EDFFXL \rf_reg<0><2>  ( .D(n952), .E(n1005), .CK(clk), .Q(\rf<0><2> ) );
  EDFFXL \rf_reg<0><1>  ( .D(n951), .E(n1005), .CK(clk), .Q(\rf<0><1> ) );
  EDFFXL \rf_reg<0><0>  ( .D(n950), .E(n1005), .CK(clk), .Q(\rf<0><0> ) );
  EDFFXL \rf_reg<10><31>  ( .D(n5), .E(n985), .CK(clk), .Q(\rf<10><31> ) );
  EDFFXL \rf_reg<10><30>  ( .D(n975), .E(n985), .CK(clk), .Q(\rf<10><30> ) );
  EDFFXL \rf_reg<10><29>  ( .D(n2), .E(n985), .CK(clk), .Q(\rf<10><29> ) );
  EDFFXL \rf_reg<10><28>  ( .D(n1), .E(n985), .CK(clk), .Q(\rf<10><28> ) );
  EDFFXL \rf_reg<10><27>  ( .D(n972), .E(n985), .CK(clk), .Q(\rf<10><27> ) );
  EDFFXL \rf_reg<10><26>  ( .D(n971), .E(n985), .CK(clk), .Q(\rf<10><26> ) );
  EDFFXL \rf_reg<10><25>  ( .D(n970), .E(n985), .CK(clk), .Q(\rf<10><25> ) );
  EDFFXL \rf_reg<10><24>  ( .D(n969), .E(n18), .CK(clk), .Q(\rf<10><24> ) );
  EDFFXL \rf_reg<10><23>  ( .D(\wd3<23> ), .E(n18), .CK(clk), .Q(\rf<10><23> )
         );
  EDFFXL \rf_reg<10><22>  ( .D(n968), .E(n18), .CK(clk), .Q(\rf<10><22> ) );
  EDFFXL \rf_reg<10><21>  ( .D(n967), .E(n18), .CK(clk), .Q(\rf<10><21> ) );
  EDFFXL \rf_reg<10><20>  ( .D(n966), .E(n985), .CK(clk), .Q(\rf<10><20> ) );
  EDFFXL \rf_reg<10><19>  ( .D(n965), .E(n985), .CK(clk), .Q(\rf<10><19> ) );
  EDFFXL \rf_reg<10><18>  ( .D(n964), .E(n985), .CK(clk), .Q(\rf<10><18> ) );
  EDFFXL \rf_reg<10><17>  ( .D(n963), .E(n985), .CK(clk), .Q(\rf<10><17> ) );
  EDFFXL \rf_reg<10><16>  ( .D(n962), .E(n985), .CK(clk), .Q(\rf<10><16> ) );
  EDFFXL \rf_reg<10><15>  ( .D(\wd3<15> ), .E(n985), .CK(clk), .Q(\rf<10><15> ) );
  EDFFXL \rf_reg<10><14>  ( .D(\wd3<14> ), .E(n985), .CK(clk), .Q(\rf<10><14> ) );
  EDFFXL \rf_reg<10><13>  ( .D(\wd3<13> ), .E(n985), .CK(clk), .Q(\rf<10><13> ) );
  EDFFXL \rf_reg<10><12>  ( .D(\wd3<12> ), .E(n985), .CK(clk), .Q(\rf<10><12> ) );
  EDFFXL \rf_reg<10><11>  ( .D(n961), .E(n985), .CK(clk), .Q(\rf<10><11> ) );
  EDFFXL \rf_reg<10><10>  ( .D(n960), .E(n985), .CK(clk), .Q(\rf<10><10> ) );
  EDFFXL \rf_reg<10><9>  ( .D(n959), .E(n985), .CK(clk), .Q(\rf<10><9> ) );
  EDFFXL \rf_reg<10><8>  ( .D(n958), .E(n985), .CK(clk), .Q(\rf<10><8> ) );
  EDFFXL \rf_reg<10><7>  ( .D(n957), .E(n18), .CK(clk), .Q(\rf<10><7> ) );
  EDFFXL \rf_reg<10><6>  ( .D(n956), .E(n18), .CK(clk), .Q(\rf<10><6> ) );
  EDFFXL \rf_reg<10><5>  ( .D(n955), .E(n18), .CK(clk), .Q(\rf<10><5> ) );
  EDFFXL \rf_reg<10><4>  ( .D(n954), .E(n18), .CK(clk), .Q(\rf<10><4> ) );
  EDFFXL \rf_reg<10><3>  ( .D(n953), .E(n18), .CK(clk), .Q(\rf<10><3> ) );
  EDFFXL \rf_reg<10><2>  ( .D(n952), .E(n18), .CK(clk), .Q(\rf<10><2> ) );
  EDFFXL \rf_reg<10><1>  ( .D(n951), .E(n18), .CK(clk), .Q(\rf<10><1> ) );
  EDFFXL \rf_reg<10><0>  ( .D(n950), .E(n18), .CK(clk), .Q(\rf<10><0> ) );
  EDFFXL \rf_reg<6><31>  ( .D(n5), .E(n993), .CK(clk), .Q(\rf<6><31> ) );
  EDFFXL \rf_reg<6><30>  ( .D(n975), .E(n993), .CK(clk), .Q(\rf<6><30> ) );
  EDFFXL \rf_reg<6><29>  ( .D(n2), .E(n993), .CK(clk), .Q(\rf<6><29> ) );
  EDFFXL \rf_reg<6><28>  ( .D(n1), .E(n993), .CK(clk), .Q(\rf<6><28> ) );
  EDFFXL \rf_reg<6><27>  ( .D(n972), .E(n993), .CK(clk), .Q(\rf<6><27> ) );
  EDFFXL \rf_reg<6><26>  ( .D(n971), .E(n993), .CK(clk), .Q(\rf<6><26> ) );
  EDFFXL \rf_reg<6><25>  ( .D(n970), .E(n993), .CK(clk), .Q(\rf<6><25> ) );
  EDFFXL \rf_reg<6><24>  ( .D(n969), .E(n16), .CK(clk), .Q(\rf<6><24> ) );
  EDFFXL \rf_reg<6><23>  ( .D(\wd3<23> ), .E(n16), .CK(clk), .Q(\rf<6><23> )
         );
  EDFFXL \rf_reg<6><22>  ( .D(n968), .E(n16), .CK(clk), .Q(\rf<6><22> ) );
  EDFFXL \rf_reg<6><21>  ( .D(n967), .E(n16), .CK(clk), .Q(\rf<6><21> ) );
  EDFFXL \rf_reg<6><20>  ( .D(n966), .E(n993), .CK(clk), .Q(\rf<6><20> ) );
  EDFFXL \rf_reg<6><19>  ( .D(n965), .E(n993), .CK(clk), .Q(\rf<6><19> ) );
  EDFFXL \rf_reg<6><18>  ( .D(n964), .E(n993), .CK(clk), .Q(\rf<6><18> ) );
  EDFFXL \rf_reg<6><17>  ( .D(n963), .E(n993), .CK(clk), .Q(\rf<6><17> ) );
  EDFFXL \rf_reg<6><16>  ( .D(n962), .E(n993), .CK(clk), .Q(\rf<6><16> ) );
  EDFFXL \rf_reg<6><15>  ( .D(\wd3<15> ), .E(n993), .CK(clk), .Q(\rf<6><15> )
         );
  EDFFXL \rf_reg<6><14>  ( .D(\wd3<14> ), .E(n993), .CK(clk), .Q(\rf<6><14> )
         );
  EDFFXL \rf_reg<6><13>  ( .D(\wd3<13> ), .E(n993), .CK(clk), .Q(\rf<6><13> )
         );
  EDFFXL \rf_reg<6><12>  ( .D(\wd3<12> ), .E(n993), .CK(clk), .Q(\rf<6><12> )
         );
  EDFFXL \rf_reg<6><11>  ( .D(n961), .E(n993), .CK(clk), .Q(\rf<6><11> ) );
  EDFFXL \rf_reg<6><10>  ( .D(n960), .E(n993), .CK(clk), .Q(\rf<6><10> ) );
  EDFFXL \rf_reg<6><9>  ( .D(n959), .E(n993), .CK(clk), .Q(\rf<6><9> ) );
  EDFFXL \rf_reg<6><8>  ( .D(n958), .E(n993), .CK(clk), .Q(\rf<6><8> ) );
  EDFFXL \rf_reg<6><7>  ( .D(n957), .E(n16), .CK(clk), .Q(\rf<6><7> ) );
  EDFFXL \rf_reg<6><6>  ( .D(n956), .E(n16), .CK(clk), .Q(\rf<6><6> ) );
  EDFFXL \rf_reg<6><5>  ( .D(n955), .E(n16), .CK(clk), .Q(\rf<6><5> ) );
  EDFFXL \rf_reg<6><4>  ( .D(n954), .E(n16), .CK(clk), .Q(\rf<6><4> ) );
  EDFFXL \rf_reg<6><3>  ( .D(n953), .E(n16), .CK(clk), .Q(\rf<6><3> ) );
  EDFFXL \rf_reg<6><2>  ( .D(n952), .E(n16), .CK(clk), .Q(\rf<6><2> ) );
  EDFFXL \rf_reg<6><1>  ( .D(n951), .E(n16), .CK(clk), .Q(\rf<6><1> ) );
  EDFFXL \rf_reg<6><0>  ( .D(n950), .E(n16), .CK(clk), .Q(\rf<6><0> ) );
  EDFFXL \rf_reg<2><31>  ( .D(n5), .E(n1001), .CK(clk), .Q(\rf<2><31> ) );
  EDFFXL \rf_reg<2><30>  ( .D(n975), .E(n1001), .CK(clk), .Q(\rf<2><30> ) );
  EDFFXL \rf_reg<2><29>  ( .D(n2), .E(n1001), .CK(clk), .Q(\rf<2><29> ) );
  EDFFXL \rf_reg<2><28>  ( .D(n1), .E(n1001), .CK(clk), .Q(\rf<2><28> ) );
  EDFFXL \rf_reg<2><27>  ( .D(n972), .E(n1001), .CK(clk), .Q(\rf<2><27> ) );
  EDFFXL \rf_reg<2><26>  ( .D(n971), .E(n1001), .CK(clk), .Q(\rf<2><26> ) );
  EDFFXL \rf_reg<2><25>  ( .D(n970), .E(n1001), .CK(clk), .Q(\rf<2><25> ) );
  EDFFXL \rf_reg<2><24>  ( .D(n969), .E(n11), .CK(clk), .Q(\rf<2><24> ) );
  EDFFXL \rf_reg<2><23>  ( .D(\wd3<23> ), .E(n11), .CK(clk), .Q(\rf<2><23> )
         );
  EDFFXL \rf_reg<2><22>  ( .D(n968), .E(n11), .CK(clk), .Q(\rf<2><22> ) );
  EDFFXL \rf_reg<2><21>  ( .D(n967), .E(n11), .CK(clk), .Q(\rf<2><21> ) );
  EDFFXL \rf_reg<2><20>  ( .D(n966), .E(n1001), .CK(clk), .Q(\rf<2><20> ) );
  EDFFXL \rf_reg<2><19>  ( .D(n965), .E(n1001), .CK(clk), .Q(\rf<2><19> ) );
  EDFFXL \rf_reg<2><18>  ( .D(n964), .E(n1001), .CK(clk), .Q(\rf<2><18> ) );
  EDFFXL \rf_reg<2><17>  ( .D(n963), .E(n1001), .CK(clk), .Q(\rf<2><17> ) );
  EDFFXL \rf_reg<2><16>  ( .D(n962), .E(n1001), .CK(clk), .Q(\rf<2><16> ) );
  EDFFXL \rf_reg<2><15>  ( .D(\wd3<15> ), .E(n1001), .CK(clk), .Q(\rf<2><15> )
         );
  EDFFXL \rf_reg<2><14>  ( .D(\wd3<14> ), .E(n1001), .CK(clk), .Q(\rf<2><14> )
         );
  EDFFXL \rf_reg<2><13>  ( .D(\wd3<13> ), .E(n1001), .CK(clk), .Q(\rf<2><13> )
         );
  EDFFXL \rf_reg<2><12>  ( .D(\wd3<12> ), .E(n1001), .CK(clk), .Q(\rf<2><12> )
         );
  EDFFXL \rf_reg<2><11>  ( .D(n961), .E(n1001), .CK(clk), .Q(\rf<2><11> ) );
  EDFFXL \rf_reg<2><10>  ( .D(n960), .E(n1001), .CK(clk), .Q(\rf<2><10> ) );
  EDFFXL \rf_reg<2><9>  ( .D(n959), .E(n1001), .CK(clk), .Q(\rf<2><9> ) );
  EDFFXL \rf_reg<2><8>  ( .D(n958), .E(n1001), .CK(clk), .Q(\rf<2><8> ) );
  EDFFXL \rf_reg<2><7>  ( .D(n957), .E(n11), .CK(clk), .Q(\rf<2><7> ) );
  EDFFXL \rf_reg<2><6>  ( .D(n956), .E(n11), .CK(clk), .Q(\rf<2><6> ) );
  EDFFXL \rf_reg<2><5>  ( .D(n955), .E(n11), .CK(clk), .Q(\rf<2><5> ) );
  EDFFXL \rf_reg<2><4>  ( .D(n954), .E(n11), .CK(clk), .Q(\rf<2><4> ) );
  EDFFXL \rf_reg<2><3>  ( .D(n953), .E(n11), .CK(clk), .Q(\rf<2><3> ) );
  EDFFXL \rf_reg<2><2>  ( .D(n952), .E(n11), .CK(clk), .Q(\rf<2><2> ) );
  EDFFXL \rf_reg<2><1>  ( .D(n951), .E(n11), .CK(clk), .Q(\rf<2><1> ) );
  EDFFXL \rf_reg<2><0>  ( .D(n950), .E(n11), .CK(clk), .Q(\rf<2><0> ) );
  EDFFXL \rf_reg<12><31>  ( .D(n5), .E(n981), .CK(clk), .Q(\rf<12><31> ) );
  EDFFXL \rf_reg<12><30>  ( .D(n975), .E(n981), .CK(clk), .Q(\rf<12><30> ) );
  EDFFXL \rf_reg<12><29>  ( .D(n2), .E(n981), .CK(clk), .Q(\rf<12><29> ) );
  EDFFXL \rf_reg<12><28>  ( .D(n1), .E(n981), .CK(clk), .Q(\rf<12><28> ) );
  EDFFXL \rf_reg<12><27>  ( .D(n972), .E(n981), .CK(clk), .Q(\rf<12><27> ) );
  EDFFXL \rf_reg<12><26>  ( .D(n971), .E(n981), .CK(clk), .Q(\rf<12><26> ) );
  EDFFXL \rf_reg<12><25>  ( .D(n970), .E(n981), .CK(clk), .Q(\rf<12><25> ) );
  EDFFXL \rf_reg<12><24>  ( .D(n969), .E(n15), .CK(clk), .Q(\rf<12><24> ) );
  EDFFXL \rf_reg<12><23>  ( .D(\wd3<23> ), .E(n15), .CK(clk), .Q(\rf<12><23> )
         );
  EDFFXL \rf_reg<12><22>  ( .D(n968), .E(n15), .CK(clk), .Q(\rf<12><22> ) );
  EDFFXL \rf_reg<12><21>  ( .D(n967), .E(n15), .CK(clk), .Q(\rf<12><21> ) );
  EDFFXL \rf_reg<12><20>  ( .D(n966), .E(n981), .CK(clk), .Q(\rf<12><20> ) );
  EDFFXL \rf_reg<12><19>  ( .D(n965), .E(n981), .CK(clk), .Q(\rf<12><19> ) );
  EDFFXL \rf_reg<12><18>  ( .D(n964), .E(n981), .CK(clk), .Q(\rf<12><18> ) );
  EDFFXL \rf_reg<12><17>  ( .D(n963), .E(n981), .CK(clk), .Q(\rf<12><17> ) );
  EDFFXL \rf_reg<12><16>  ( .D(n962), .E(n981), .CK(clk), .Q(\rf<12><16> ) );
  EDFFXL \rf_reg<12><15>  ( .D(\wd3<15> ), .E(n981), .CK(clk), .Q(\rf<12><15> ) );
  EDFFXL \rf_reg<12><14>  ( .D(\wd3<14> ), .E(n981), .CK(clk), .Q(\rf<12><14> ) );
  EDFFXL \rf_reg<12><13>  ( .D(\wd3<13> ), .E(n981), .CK(clk), .Q(\rf<12><13> ) );
  EDFFXL \rf_reg<12><12>  ( .D(\wd3<12> ), .E(n981), .CK(clk), .Q(\rf<12><12> ) );
  EDFFXL \rf_reg<12><11>  ( .D(n961), .E(n981), .CK(clk), .Q(\rf<12><11> ) );
  EDFFXL \rf_reg<12><10>  ( .D(n960), .E(n981), .CK(clk), .Q(\rf<12><10> ) );
  EDFFXL \rf_reg<12><9>  ( .D(n959), .E(n981), .CK(clk), .Q(\rf<12><9> ) );
  EDFFXL \rf_reg<12><8>  ( .D(n958), .E(n981), .CK(clk), .Q(\rf<12><8> ) );
  EDFFXL \rf_reg<12><7>  ( .D(n957), .E(n15), .CK(clk), .Q(\rf<12><7> ) );
  EDFFXL \rf_reg<12><6>  ( .D(n956), .E(n15), .CK(clk), .Q(\rf<12><6> ) );
  EDFFXL \rf_reg<12><5>  ( .D(n955), .E(n15), .CK(clk), .Q(\rf<12><5> ) );
  EDFFXL \rf_reg<12><4>  ( .D(n954), .E(n15), .CK(clk), .Q(\rf<12><4> ) );
  EDFFXL \rf_reg<12><3>  ( .D(n953), .E(n15), .CK(clk), .Q(\rf<12><3> ) );
  EDFFXL \rf_reg<12><2>  ( .D(n952), .E(n15), .CK(clk), .Q(\rf<12><2> ) );
  EDFFXL \rf_reg<12><1>  ( .D(n951), .E(n15), .CK(clk), .Q(\rf<12><1> ) );
  EDFFXL \rf_reg<12><0>  ( .D(n950), .E(n15), .CK(clk), .Q(\rf<12><0> ) );
  BUFX20 U4 ( .A(n973), .Y(n1) );
  BUFX1 U5 ( .A(\wd3<28> ), .Y(n973) );
  BUFX8 U6 ( .A(\wd3<27> ), .Y(n972) );
  BUFX20 U7 ( .A(\wd3<30> ), .Y(n975) );
  BUFX20 U8 ( .A(n974), .Y(n2) );
  BUFX1 U9 ( .A(\wd3<29> ), .Y(n974) );
  BUFX20 U10 ( .A(\wd3<31> ), .Y(n5) );
  OAI2BB2X1 U11 ( .B0(n1017), .B1(n1007), .A0N(N503), .A1N(n1007), .Y(
        \rd1<31> ) );
  OAI2BB2X1 U12 ( .B0(n1010), .B1(n1017), .A0N(N536), .A1N(n1010), .Y(
        \rd2<31> ) );
  AND4X2 U13 ( .A(N15), .B(N14), .C(N13), .D(N12), .Y(n3) );
  AND4X2 U14 ( .A(N19), .B(N18), .C(N17), .D(n944), .Y(n4) );
  INVX12 U15 ( .A(\r15<31> ), .Y(n1017) );
  CLKINVX3 U16 ( .A(n936), .Y(n944) );
  CLKINVX3 U17 ( .A(n780), .Y(n786) );
  CLKINVX3 U18 ( .A(n780), .Y(n785) );
  CLKINVX3 U19 ( .A(n788), .Y(n784) );
  CLKINVX3 U20 ( .A(n788), .Y(n783) );
  CLKINVX3 U21 ( .A(n779), .Y(n782) );
  CLKINVX3 U22 ( .A(n779), .Y(n781) );
  CLKINVX3 U23 ( .A(n779), .Y(n787) );
  CLKINVX3 U24 ( .A(n938), .Y(n949) );
  CLKINVX3 U25 ( .A(n936), .Y(n948) );
  CLKINVX3 U26 ( .A(n939), .Y(n947) );
  CLKINVX3 U27 ( .A(n936), .Y(n946) );
  CLKINVX3 U28 ( .A(n936), .Y(n945) );
  CLKINVX3 U29 ( .A(n940), .Y(n943) );
  INVX1 U30 ( .A(n773), .Y(n780) );
  INVX1 U31 ( .A(n773), .Y(n779) );
  INVX1 U32 ( .A(n774), .Y(n775) );
  INVX1 U33 ( .A(n774), .Y(n776) );
  INVX1 U34 ( .A(n774), .Y(n777) );
  INVX1 U35 ( .A(n773), .Y(n778) );
  INVX1 U36 ( .A(n937), .Y(n938) );
  INVX1 U37 ( .A(n937), .Y(n939) );
  INVX1 U38 ( .A(N16), .Y(n940) );
  INVX1 U39 ( .A(N16), .Y(n941) );
  INVX1 U40 ( .A(n937), .Y(n942) );
  CLKINVX3 U41 ( .A(n1015), .Y(n765) );
  CLKINVX3 U42 ( .A(n1015), .Y(n766) );
  CLKINVX3 U43 ( .A(n1013), .Y(n929) );
  CLKINVX3 U44 ( .A(n1013), .Y(n930) );
  CLKINVX3 U45 ( .A(n764), .Y(n771) );
  CLKINVX3 U46 ( .A(n764), .Y(n770) );
  CLKINVX3 U47 ( .A(n764), .Y(n769) );
  CLKINVX3 U48 ( .A(n764), .Y(n768) );
  CLKINVX3 U49 ( .A(n1015), .Y(n767) );
  CLKINVX3 U50 ( .A(n1013), .Y(n935) );
  CLKINVX3 U51 ( .A(n1013), .Y(n934) );
  CLKINVX3 U52 ( .A(n928), .Y(n933) );
  CLKINVX3 U53 ( .A(n928), .Y(n932) );
  CLKINVX3 U54 ( .A(n1013), .Y(n931) );
  INVX1 U55 ( .A(n778), .Y(n774) );
  INVX1 U56 ( .A(n788), .Y(n773) );
  INVX1 U57 ( .A(n936), .Y(n937) );
  CLKINVX3 U58 ( .A(n1016), .Y(n759) );
  CLKINVX3 U59 ( .A(n1014), .Y(n923) );
  CLKINVX3 U60 ( .A(n3), .Y(n1009) );
  CLKINVX3 U61 ( .A(n4), .Y(n1012) );
  CLKINVX3 U62 ( .A(n4), .Y(n1011) );
  CLKINVX3 U63 ( .A(n3), .Y(n1008) );
  CLKINVX3 U64 ( .A(n761), .Y(n762) );
  CLKINVX3 U65 ( .A(n925), .Y(n926) );
  INVX1 U66 ( .A(N16), .Y(n936) );
  INVX1 U67 ( .A(n772), .Y(n764) );
  INVX1 U68 ( .A(n930), .Y(n928) );
  CLKINVX3 U69 ( .A(n4), .Y(n1010) );
  CLKINVX3 U70 ( .A(n3), .Y(n1007) );
  CLKINVX3 U71 ( .A(n761), .Y(n763) );
  INVX1 U72 ( .A(N14), .Y(n761) );
  CLKINVX3 U73 ( .A(n925), .Y(n927) );
  INVX1 U74 ( .A(N18), .Y(n925) );
  INVX1 U75 ( .A(n1015), .Y(n772) );
  CLKINVX3 U76 ( .A(n1016), .Y(n760) );
  CLKINVX3 U77 ( .A(n1014), .Y(n924) );
  CLKINVX3 U78 ( .A(n1004), .Y(n1003) );
  CLKINVX3 U79 ( .A(n1002), .Y(n1001) );
  CLKINVX3 U80 ( .A(n1000), .Y(n999) );
  CLKINVX3 U81 ( .A(n998), .Y(n997) );
  CLKINVX3 U82 ( .A(n996), .Y(n995) );
  CLKINVX3 U83 ( .A(n994), .Y(n993) );
  CLKINVX3 U84 ( .A(n992), .Y(n991) );
  CLKINVX3 U85 ( .A(n990), .Y(n989) );
  CLKINVX3 U86 ( .A(n988), .Y(n987) );
  CLKINVX3 U87 ( .A(n986), .Y(n985) );
  CLKINVX3 U88 ( .A(n984), .Y(n983) );
  CLKINVX3 U89 ( .A(n982), .Y(n981) );
  CLKINVX3 U90 ( .A(n980), .Y(n979) );
  CLKINVX3 U91 ( .A(n978), .Y(n977) );
  CLKINVX3 U92 ( .A(n1006), .Y(n1005) );
  INVX1 U93 ( .A(N12), .Y(n788) );
  INVX1 U94 ( .A(n9), .Y(n1006) );
  INVX1 U95 ( .A(n7), .Y(n988) );
  INVX1 U96 ( .A(n8), .Y(n980) );
  INVX1 U97 ( .A(n10), .Y(n1004) );
  INVX1 U98 ( .A(n13), .Y(n998) );
  INVX1 U99 ( .A(n6), .Y(n996) );
  INVX1 U100 ( .A(n16), .Y(n994) );
  INVX1 U101 ( .A(n17), .Y(n992) );
  INVX1 U102 ( .A(n11), .Y(n1002) );
  INVX1 U103 ( .A(n12), .Y(n1000) );
  INVX1 U104 ( .A(n14), .Y(n990) );
  INVX1 U105 ( .A(n15), .Y(n982) );
  INVX1 U106 ( .A(n18), .Y(n986) );
  INVX1 U107 ( .A(n20), .Y(n984) );
  INVX1 U108 ( .A(n19), .Y(n978) );
  INVX1 U109 ( .A(\r15<26> ), .Y(n1022) );
  INVX1 U110 ( .A(\r15<27> ), .Y(n1021) );
  INVX1 U111 ( .A(\r15<28> ), .Y(n1020) );
  INVX1 U112 ( .A(\r15<29> ), .Y(n1019) );
  INVX1 U113 ( .A(\r15<30> ), .Y(n1018) );
  BUFX3 U114 ( .A(\wd3<26> ), .Y(n971) );
  INVX1 U115 ( .A(\r15<21> ), .Y(n1027) );
  INVX1 U116 ( .A(\r15<22> ), .Y(n1026) );
  INVX1 U117 ( .A(\r15<23> ), .Y(n1025) );
  INVX1 U118 ( .A(\r15<24> ), .Y(n1024) );
  INVX1 U119 ( .A(\r15<25> ), .Y(n1023) );
  BUFX3 U120 ( .A(\wd3<21> ), .Y(n967) );
  BUFX3 U121 ( .A(\wd3<22> ), .Y(n968) );
  BUFX3 U122 ( .A(\wd3<24> ), .Y(n969) );
  BUFX3 U123 ( .A(\wd3<25> ), .Y(n970) );
  INVX1 U124 ( .A(\r15<16> ), .Y(n1032) );
  INVX1 U125 ( .A(\r15<17> ), .Y(n1031) );
  INVX1 U126 ( .A(\r15<18> ), .Y(n1030) );
  INVX1 U127 ( .A(\r15<19> ), .Y(n1029) );
  INVX1 U128 ( .A(\r15<20> ), .Y(n1028) );
  BUFX3 U129 ( .A(\wd3<16> ), .Y(n962) );
  BUFX3 U130 ( .A(\wd3<17> ), .Y(n963) );
  BUFX3 U131 ( .A(\wd3<18> ), .Y(n964) );
  BUFX3 U132 ( .A(\wd3<19> ), .Y(n965) );
  BUFX3 U133 ( .A(\wd3<20> ), .Y(n966) );
  INVX1 U134 ( .A(\r15<11> ), .Y(n1037) );
  INVX1 U135 ( .A(\r15<12> ), .Y(n1036) );
  INVX1 U136 ( .A(\r15<13> ), .Y(n1035) );
  INVX1 U137 ( .A(\r15<14> ), .Y(n1034) );
  INVX1 U138 ( .A(\r15<15> ), .Y(n1033) );
  BUFX3 U139 ( .A(\wd3<10> ), .Y(n960) );
  BUFX3 U140 ( .A(\wd3<11> ), .Y(n961) );
  INVX1 U141 ( .A(\r15<9> ), .Y(n1039) );
  INVX1 U142 ( .A(\r15<6> ), .Y(n1042) );
  INVX1 U143 ( .A(\r15<7> ), .Y(n1041) );
  INVX1 U144 ( .A(\r15<8> ), .Y(n1040) );
  INVX1 U145 ( .A(\r15<10> ), .Y(n1038) );
  BUFX3 U146 ( .A(\wd3<5> ), .Y(n955) );
  BUFX3 U147 ( .A(\wd3<6> ), .Y(n956) );
  BUFX3 U148 ( .A(\wd3<7> ), .Y(n957) );
  BUFX3 U149 ( .A(\wd3<8> ), .Y(n958) );
  BUFX3 U150 ( .A(\wd3<9> ), .Y(n959) );
  INVX1 U151 ( .A(\r15<1> ), .Y(n1047) );
  INVX1 U152 ( .A(\r15<2> ), .Y(n1046) );
  INVX1 U153 ( .A(\r15<3> ), .Y(n1045) );
  INVX1 U154 ( .A(\r15<4> ), .Y(n1044) );
  INVX1 U155 ( .A(\r15<5> ), .Y(n1043) );
  BUFX3 U156 ( .A(\wd3<1> ), .Y(n951) );
  BUFX3 U157 ( .A(\wd3<2> ), .Y(n952) );
  BUFX3 U158 ( .A(\wd3<3> ), .Y(n953) );
  BUFX3 U159 ( .A(\wd3<4> ), .Y(n954) );
  INVX1 U160 ( .A(\r15<0> ), .Y(n1048) );
  BUFX3 U161 ( .A(\wd3<0> ), .Y(n950) );
  INVX1 U162 ( .A(N19), .Y(n1014) );
  INVX1 U163 ( .A(N13), .Y(n1015) );
  INVX1 U164 ( .A(N17), .Y(n1013) );
  INVX1 U165 ( .A(N15), .Y(n1016) );
  AND3X2 U166 ( .A(n537), .B(n976), .C(n543), .Y(n6) );
  AND3X2 U167 ( .A(n537), .B(n976), .C(n548), .Y(n7) );
  AND3X2 U168 ( .A(n537), .B(n976), .C(n553), .Y(n8) );
  AND3X2 U169 ( .A(n534), .B(n535), .C(n976), .Y(n9) );
  AND3X2 U170 ( .A(n976), .B(n534), .C(n537), .Y(n10) );
  AND3X2 U171 ( .A(n976), .B(n534), .C(n539), .Y(n11) );
  AND3X2 U172 ( .A(n976), .B(n534), .C(n541), .Y(n12) );
  AND3X2 U173 ( .A(n976), .B(n535), .C(n543), .Y(n13) );
  AND3X2 U174 ( .A(n976), .B(n535), .C(n548), .Y(n14) );
  AND3X2 U175 ( .A(n976), .B(n535), .C(n553), .Y(n15) );
  AND3X2 U176 ( .A(n539), .B(n976), .C(n543), .Y(n16) );
  AND3X2 U177 ( .A(n541), .B(n976), .C(n543), .Y(n17) );
  AND3X2 U178 ( .A(n539), .B(n976), .C(n548), .Y(n18) );
  AND3X2 U179 ( .A(n539), .B(n976), .C(n553), .Y(n19) );
  AND3X2 U180 ( .A(n541), .B(n976), .C(n548), .Y(n20) );
  MX4X1 U181 ( .A(n922), .B(n920), .C(n921), .D(n919), .S0(n924), .S1(n927), 
        .Y(N536) );
  MX4X1 U182 ( .A(\rf<0><31> ), .B(\rf<1><31> ), .C(\rf<2><31> ), .D(
        \rf<3><31> ), .S0(n945), .S1(N17), .Y(n922) );
  MX4X1 U183 ( .A(\rf<8><31> ), .B(\rf<9><31> ), .C(\rf<10><31> ), .D(
        \rf<11><31> ), .S0(n945), .S1(n931), .Y(n920) );
  MX4X1 U184 ( .A(n758), .B(n756), .C(n757), .D(n755), .S0(n760), .S1(n763), 
        .Y(N503) );
  MX4X1 U185 ( .A(\rf<0><31> ), .B(\rf<1><31> ), .C(\rf<2><31> ), .D(
        \rf<3><31> ), .S0(n787), .S1(n767), .Y(n758) );
  MX4X1 U186 ( .A(\rf<8><31> ), .B(\rf<9><31> ), .C(\rf<10><31> ), .D(
        \rf<11><31> ), .S0(n774), .S1(n767), .Y(n756) );
  OAI2BB2X1 U187 ( .B0(n1011), .B1(n1022), .A0N(N541), .A1N(n1012), .Y(
        \rd2<26> ) );
  MX4X1 U188 ( .A(n898), .B(n896), .C(n897), .D(n895), .S0(n924), .S1(n927), 
        .Y(N541) );
  MX4X1 U189 ( .A(\rf<0><26> ), .B(\rf<1><26> ), .C(\rf<2><26> ), .D(
        \rf<3><26> ), .S0(n946), .S1(n932), .Y(n898) );
  MX4X1 U190 ( .A(\rf<8><26> ), .B(\rf<9><26> ), .C(\rf<10><26> ), .D(
        \rf<11><26> ), .S0(n946), .S1(n932), .Y(n896) );
  OAI2BB2X1 U191 ( .B0(n1010), .B1(n1021), .A0N(N540), .A1N(n1012), .Y(
        \rd2<27> ) );
  MX4X1 U192 ( .A(n902), .B(n900), .C(n901), .D(n899), .S0(n924), .S1(n927), 
        .Y(N540) );
  MX4X1 U193 ( .A(\rf<0><27> ), .B(\rf<1><27> ), .C(\rf<2><27> ), .D(
        \rf<3><27> ), .S0(n946), .S1(n932), .Y(n902) );
  MX4X1 U194 ( .A(\rf<8><27> ), .B(\rf<9><27> ), .C(\rf<10><27> ), .D(
        \rf<11><27> ), .S0(n946), .S1(n932), .Y(n900) );
  OAI2BB2X1 U195 ( .B0(n1010), .B1(n1020), .A0N(N539), .A1N(n1012), .Y(
        \rd2<28> ) );
  MX4X1 U196 ( .A(n906), .B(n904), .C(n905), .D(n903), .S0(n924), .S1(n927), 
        .Y(N539) );
  MX4X1 U197 ( .A(\rf<0><28> ), .B(\rf<1><28> ), .C(\rf<2><28> ), .D(
        \rf<3><28> ), .S0(n945), .S1(n931), .Y(n906) );
  MX4X1 U198 ( .A(\rf<8><28> ), .B(\rf<9><28> ), .C(\rf<10><28> ), .D(
        \rf<11><28> ), .S0(n945), .S1(n931), .Y(n904) );
  OAI2BB2X1 U199 ( .B0(n1010), .B1(n1019), .A0N(N538), .A1N(n1012), .Y(
        \rd2<29> ) );
  MX4X1 U200 ( .A(n912), .B(n910), .C(n911), .D(n909), .S0(n924), .S1(n927), 
        .Y(N538) );
  MX2X1 U201 ( .A(n907), .B(n908), .S0(n932), .Y(n909) );
  MX4X1 U202 ( .A(\rf<0><29> ), .B(\rf<1><29> ), .C(\rf<2><29> ), .D(
        \rf<3><29> ), .S0(n945), .S1(n931), .Y(n912) );
  OAI2BB2X1 U203 ( .B0(n1010), .B1(n1018), .A0N(N537), .A1N(n1012), .Y(
        \rd2<30> ) );
  MX4X1 U204 ( .A(n918), .B(n916), .C(n917), .D(n915), .S0(n924), .S1(n927), 
        .Y(N537) );
  MX2X1 U205 ( .A(n913), .B(n914), .S0(n929), .Y(n915) );
  MX4X1 U206 ( .A(\rf<0><30> ), .B(\rf<1><30> ), .C(\rf<2><30> ), .D(
        \rf<3><30> ), .S0(n945), .S1(n931), .Y(n918) );
  OAI2BB2X1 U207 ( .B0(n1022), .B1(n1008), .A0N(N508), .A1N(n1009), .Y(
        \rd1<26> ) );
  MX4X1 U208 ( .A(n734), .B(n732), .C(n733), .D(n731), .S0(n760), .S1(n763), 
        .Y(N508) );
  MX4X1 U209 ( .A(\rf<0><26> ), .B(\rf<1><26> ), .C(\rf<2><26> ), .D(
        \rf<3><26> ), .S0(n781), .S1(n772), .Y(n734) );
  MX4X1 U210 ( .A(\rf<8><26> ), .B(\rf<9><26> ), .C(\rf<10><26> ), .D(
        \rf<11><26> ), .S0(n781), .S1(n767), .Y(n732) );
  OAI2BB2X1 U211 ( .B0(n1021), .B1(n1007), .A0N(N507), .A1N(n1009), .Y(
        \rd1<27> ) );
  MX4X1 U212 ( .A(n738), .B(n736), .C(n737), .D(n735), .S0(n760), .S1(n763), 
        .Y(N507) );
  MX4X1 U213 ( .A(\rf<0><27> ), .B(\rf<1><27> ), .C(\rf<2><27> ), .D(
        \rf<3><27> ), .S0(n781), .S1(n767), .Y(n738) );
  MX4X1 U214 ( .A(\rf<8><27> ), .B(\rf<9><27> ), .C(\rf<10><27> ), .D(
        \rf<11><27> ), .S0(n781), .S1(n766), .Y(n736) );
  OAI2BB2X1 U215 ( .B0(n1020), .B1(n1007), .A0N(N506), .A1N(n1009), .Y(
        \rd1<28> ) );
  MX4X1 U216 ( .A(n742), .B(n740), .C(n741), .D(n739), .S0(n760), .S1(n763), 
        .Y(N506) );
  MX4X1 U217 ( .A(\rf<0><28> ), .B(\rf<1><28> ), .C(\rf<2><28> ), .D(
        \rf<3><28> ), .S0(n783), .S1(n767), .Y(n742) );
  MX4X1 U218 ( .A(\rf<8><28> ), .B(\rf<9><28> ), .C(\rf<10><28> ), .D(
        \rf<11><28> ), .S0(n783), .S1(n767), .Y(n740) );
  OAI2BB2X1 U219 ( .B0(n1019), .B1(n1007), .A0N(N505), .A1N(n1009), .Y(
        \rd1<29> ) );
  MX4X1 U220 ( .A(n748), .B(n746), .C(n747), .D(n745), .S0(n760), .S1(n763), 
        .Y(N505) );
  MX2X1 U221 ( .A(n743), .B(n744), .S0(n768), .Y(n745) );
  MX4X1 U222 ( .A(\rf<0><29> ), .B(\rf<1><29> ), .C(\rf<2><29> ), .D(
        \rf<3><29> ), .S0(n784), .S1(n767), .Y(n748) );
  OAI2BB2X1 U223 ( .B0(n1018), .B1(n1007), .A0N(N504), .A1N(n1009), .Y(
        \rd1<30> ) );
  MX4X1 U224 ( .A(n754), .B(n752), .C(n753), .D(n751), .S0(n760), .S1(n763), 
        .Y(N504) );
  MX2X1 U225 ( .A(n749), .B(n750), .S0(n769), .Y(n751) );
  MX4X1 U226 ( .A(\rf<0><30> ), .B(\rf<1><30> ), .C(\rf<2><30> ), .D(
        \rf<3><30> ), .S0(n787), .S1(n767), .Y(n754) );
  OAI2BB2X1 U227 ( .B0(n1011), .B1(n1027), .A0N(N546), .A1N(n1011), .Y(
        \rd2<21> ) );
  MX4X1 U228 ( .A(n878), .B(n876), .C(n877), .D(n875), .S0(n924), .S1(n927), 
        .Y(N546) );
  MX4X1 U229 ( .A(\rf<0><21> ), .B(\rf<1><21> ), .C(\rf<2><21> ), .D(
        \rf<3><21> ), .S0(n948), .S1(n934), .Y(n878) );
  MX4X1 U230 ( .A(\rf<8><21> ), .B(\rf<9><21> ), .C(\rf<10><21> ), .D(
        \rf<11><21> ), .S0(n948), .S1(n934), .Y(n876) );
  OAI2BB2X1 U231 ( .B0(n1011), .B1(n1026), .A0N(N545), .A1N(n1010), .Y(
        \rd2<22> ) );
  MX4X1 U232 ( .A(n882), .B(n880), .C(n881), .D(n879), .S0(n924), .S1(n927), 
        .Y(N545) );
  MX4X1 U233 ( .A(\rf<0><22> ), .B(\rf<1><22> ), .C(\rf<2><22> ), .D(
        \rf<3><22> ), .S0(n947), .S1(n933), .Y(n882) );
  MX4X1 U234 ( .A(\rf<8><22> ), .B(\rf<9><22> ), .C(\rf<10><22> ), .D(
        \rf<11><22> ), .S0(n947), .S1(n933), .Y(n880) );
  OAI2BB2X1 U235 ( .B0(n1011), .B1(n1025), .A0N(N544), .A1N(n1012), .Y(
        \rd2<23> ) );
  MX4X1 U236 ( .A(n886), .B(n884), .C(n885), .D(n883), .S0(n924), .S1(n927), 
        .Y(N544) );
  MX4X1 U237 ( .A(\rf<0><23> ), .B(\rf<1><23> ), .C(\rf<2><23> ), .D(
        \rf<3><23> ), .S0(n947), .S1(n933), .Y(n886) );
  MX4X1 U238 ( .A(\rf<8><23> ), .B(\rf<9><23> ), .C(\rf<10><23> ), .D(
        \rf<11><23> ), .S0(n947), .S1(n933), .Y(n884) );
  OAI2BB2X1 U239 ( .B0(n1011), .B1(n1024), .A0N(N543), .A1N(n1012), .Y(
        \rd2<24> ) );
  MX4X1 U240 ( .A(n890), .B(n888), .C(n889), .D(n887), .S0(n924), .S1(n927), 
        .Y(N543) );
  MX4X1 U241 ( .A(\rf<0><24> ), .B(\rf<1><24> ), .C(\rf<2><24> ), .D(
        \rf<3><24> ), .S0(n947), .S1(n933), .Y(n890) );
  MX4X1 U242 ( .A(\rf<8><24> ), .B(\rf<9><24> ), .C(\rf<10><24> ), .D(
        \rf<11><24> ), .S0(n947), .S1(n933), .Y(n888) );
  OAI2BB2X1 U243 ( .B0(n1011), .B1(n1023), .A0N(N542), .A1N(n1012), .Y(
        \rd2<25> ) );
  MX4X1 U244 ( .A(n894), .B(n892), .C(n893), .D(n891), .S0(n924), .S1(n927), 
        .Y(N542) );
  MX4X1 U245 ( .A(\rf<0><25> ), .B(\rf<1><25> ), .C(\rf<2><25> ), .D(
        \rf<3><25> ), .S0(n946), .S1(n932), .Y(n894) );
  MX4X1 U246 ( .A(\rf<8><25> ), .B(\rf<9><25> ), .C(\rf<10><25> ), .D(
        \rf<11><25> ), .S0(n946), .S1(n932), .Y(n892) );
  OAI2BB2X1 U247 ( .B0(n1027), .B1(n1008), .A0N(N513), .A1N(n1008), .Y(
        \rd1<21> ) );
  MX4X1 U248 ( .A(n714), .B(n712), .C(n713), .D(n711), .S0(n760), .S1(n763), 
        .Y(N513) );
  MX4X1 U249 ( .A(\rf<0><21> ), .B(\rf<1><21> ), .C(\rf<2><21> ), .D(
        \rf<3><21> ), .S0(n783), .S1(n768), .Y(n714) );
  MX4X1 U250 ( .A(\rf<8><21> ), .B(\rf<9><21> ), .C(\rf<10><21> ), .D(
        \rf<11><21> ), .S0(n783), .S1(n768), .Y(n712) );
  OAI2BB2X1 U251 ( .B0(n1026), .B1(n1008), .A0N(N512), .A1N(n1007), .Y(
        \rd1<22> ) );
  MX4X1 U252 ( .A(n718), .B(n716), .C(n717), .D(n715), .S0(n760), .S1(n763), 
        .Y(N512) );
  MX4X1 U253 ( .A(\rf<0><22> ), .B(\rf<1><22> ), .C(\rf<2><22> ), .D(
        \rf<3><22> ), .S0(n782), .S1(n769), .Y(n718) );
  MX4X1 U254 ( .A(\rf<8><22> ), .B(\rf<9><22> ), .C(\rf<10><22> ), .D(
        \rf<11><22> ), .S0(n782), .S1(n769), .Y(n716) );
  OAI2BB2X1 U255 ( .B0(n1025), .B1(n1008), .A0N(N511), .A1N(n1009), .Y(
        \rd1<23> ) );
  MX4X1 U256 ( .A(n722), .B(n720), .C(n721), .D(n719), .S0(n760), .S1(n763), 
        .Y(N511) );
  MX4X1 U257 ( .A(\rf<0><23> ), .B(\rf<1><23> ), .C(\rf<2><23> ), .D(
        \rf<3><23> ), .S0(n782), .S1(n771), .Y(n722) );
  MX4X1 U258 ( .A(\rf<8><23> ), .B(\rf<9><23> ), .C(\rf<10><23> ), .D(
        \rf<11><23> ), .S0(n782), .S1(n771), .Y(n720) );
  OAI2BB2X1 U259 ( .B0(n1024), .B1(n1008), .A0N(N510), .A1N(n1009), .Y(
        \rd1<24> ) );
  MX4X1 U260 ( .A(n726), .B(n724), .C(n725), .D(n723), .S0(n760), .S1(n763), 
        .Y(N510) );
  MX4X1 U261 ( .A(\rf<0><24> ), .B(\rf<1><24> ), .C(\rf<2><24> ), .D(
        \rf<3><24> ), .S0(n782), .S1(n770), .Y(n726) );
  MX4X1 U262 ( .A(\rf<8><24> ), .B(\rf<9><24> ), .C(\rf<10><24> ), .D(
        \rf<11><24> ), .S0(n782), .S1(n770), .Y(n724) );
  OAI2BB2X1 U263 ( .B0(n1023), .B1(n1008), .A0N(N509), .A1N(n1009), .Y(
        \rd1<25> ) );
  MX4X1 U264 ( .A(n730), .B(n728), .C(n729), .D(n727), .S0(n760), .S1(n763), 
        .Y(N509) );
  MX4X1 U265 ( .A(\rf<0><25> ), .B(\rf<1><25> ), .C(\rf<2><25> ), .D(
        \rf<3><25> ), .S0(n781), .S1(n766), .Y(n730) );
  MX4X1 U266 ( .A(\rf<8><25> ), .B(\rf<9><25> ), .C(\rf<10><25> ), .D(
        \rf<11><25> ), .S0(n781), .S1(n766), .Y(n728) );
  OAI2BB2X1 U267 ( .B0(n1011), .B1(n1032), .A0N(N551), .A1N(n1012), .Y(
        \rd2<16> ) );
  MX4X1 U268 ( .A(n858), .B(n856), .C(n857), .D(n855), .S0(n923), .S1(n926), 
        .Y(N551) );
  MX4X1 U269 ( .A(\rf<0><16> ), .B(\rf<1><16> ), .C(\rf<2><16> ), .D(
        \rf<3><16> ), .S0(n949), .S1(n933), .Y(n858) );
  MX4X1 U270 ( .A(\rf<8><16> ), .B(\rf<9><16> ), .C(\rf<10><16> ), .D(
        \rf<11><16> ), .S0(n949), .S1(n935), .Y(n856) );
  OAI2BB2X1 U271 ( .B0(n1011), .B1(n1031), .A0N(N550), .A1N(n1011), .Y(
        \rd2<17> ) );
  MX4X1 U272 ( .A(n862), .B(n860), .C(n861), .D(n859), .S0(n923), .S1(n926), 
        .Y(N550) );
  MX4X1 U273 ( .A(\rf<0><17> ), .B(\rf<1><17> ), .C(\rf<2><17> ), .D(
        \rf<3><17> ), .S0(n949), .S1(n932), .Y(n862) );
  MX4X1 U274 ( .A(\rf<8><17> ), .B(\rf<9><17> ), .C(\rf<10><17> ), .D(
        \rf<11><17> ), .S0(n949), .S1(n934), .Y(n860) );
  OAI2BB2X1 U275 ( .B0(n1011), .B1(n1030), .A0N(N549), .A1N(n1012), .Y(
        \rd2<18> ) );
  MX4X1 U276 ( .A(n866), .B(n864), .C(n865), .D(n863), .S0(n923), .S1(n926), 
        .Y(N549) );
  MX4X1 U277 ( .A(\rf<0><18> ), .B(\rf<1><18> ), .C(\rf<2><18> ), .D(
        \rf<3><18> ), .S0(n949), .S1(n935), .Y(n866) );
  MX4X1 U278 ( .A(\rf<8><18> ), .B(\rf<9><18> ), .C(\rf<10><18> ), .D(
        \rf<11><18> ), .S0(n949), .S1(n933), .Y(n864) );
  OAI2BB2X1 U279 ( .B0(n1011), .B1(n1029), .A0N(N548), .A1N(n1012), .Y(
        \rd2<19> ) );
  MX4X1 U280 ( .A(n870), .B(n868), .C(n869), .D(n867), .S0(n923), .S1(n926), 
        .Y(N548) );
  MX4X1 U281 ( .A(\rf<0><19> ), .B(\rf<1><19> ), .C(\rf<2><19> ), .D(
        \rf<3><19> ), .S0(n948), .S1(n934), .Y(n870) );
  MX4X1 U282 ( .A(\rf<8><19> ), .B(\rf<9><19> ), .C(\rf<10><19> ), .D(
        \rf<11><19> ), .S0(n948), .S1(n934), .Y(n868) );
  OAI2BB2X1 U283 ( .B0(n1011), .B1(n1028), .A0N(N547), .A1N(n1012), .Y(
        \rd2<20> ) );
  MX4X1 U284 ( .A(n874), .B(n872), .C(n873), .D(n871), .S0(n924), .S1(n927), 
        .Y(N547) );
  MX4X1 U285 ( .A(\rf<0><20> ), .B(\rf<1><20> ), .C(\rf<2><20> ), .D(
        \rf<3><20> ), .S0(n948), .S1(n934), .Y(n874) );
  MX4X1 U286 ( .A(\rf<8><20> ), .B(\rf<9><20> ), .C(\rf<10><20> ), .D(
        \rf<11><20> ), .S0(n948), .S1(n934), .Y(n872) );
  OAI2BB2X1 U287 ( .B0(n1032), .B1(n1008), .A0N(N518), .A1N(n1009), .Y(
        \rd1<16> ) );
  MX4X1 U288 ( .A(n694), .B(n692), .C(n693), .D(n691), .S0(n759), .S1(n762), 
        .Y(N518) );
  MX4X1 U289 ( .A(\rf<0><16> ), .B(\rf<1><16> ), .C(\rf<2><16> ), .D(
        \rf<3><16> ), .S0(n784), .S1(n769), .Y(n694) );
  MX4X1 U290 ( .A(\rf<8><16> ), .B(\rf<9><16> ), .C(\rf<10><16> ), .D(
        \rf<11><16> ), .S0(n784), .S1(n769), .Y(n692) );
  OAI2BB2X1 U291 ( .B0(n1031), .B1(n1007), .A0N(N517), .A1N(n1008), .Y(
        \rd1<17> ) );
  MX4X1 U292 ( .A(n698), .B(n696), .C(n697), .D(n695), .S0(n759), .S1(n762), 
        .Y(N517) );
  MX4X1 U293 ( .A(\rf<0><17> ), .B(\rf<1><17> ), .C(\rf<2><17> ), .D(
        \rf<3><17> ), .S0(n784), .S1(n769), .Y(n698) );
  MX4X1 U294 ( .A(\rf<8><17> ), .B(\rf<9><17> ), .C(\rf<10><17> ), .D(
        \rf<11><17> ), .S0(n784), .S1(n769), .Y(n696) );
  OAI2BB2X1 U295 ( .B0(n1030), .B1(n1008), .A0N(N516), .A1N(n1009), .Y(
        \rd1<18> ) );
  MX4X1 U296 ( .A(n702), .B(n700), .C(n701), .D(n699), .S0(n759), .S1(n762), 
        .Y(N516) );
  MX4X1 U297 ( .A(\rf<0><18> ), .B(\rf<1><18> ), .C(\rf<2><18> ), .D(
        \rf<3><18> ), .S0(n784), .S1(n769), .Y(n702) );
  MX4X1 U298 ( .A(\rf<8><18> ), .B(\rf<9><18> ), .C(\rf<10><18> ), .D(
        \rf<11><18> ), .S0(n784), .S1(n769), .Y(n700) );
  OAI2BB2X1 U299 ( .B0(n1029), .B1(n1008), .A0N(N515), .A1N(n1008), .Y(
        \rd1<19> ) );
  MX4X1 U300 ( .A(n706), .B(n704), .C(n705), .D(n703), .S0(n759), .S1(n762), 
        .Y(N515) );
  MX4X1 U301 ( .A(\rf<0><19> ), .B(\rf<1><19> ), .C(\rf<2><19> ), .D(
        \rf<3><19> ), .S0(n783), .S1(n768), .Y(n706) );
  MX4X1 U302 ( .A(\rf<8><19> ), .B(\rf<9><19> ), .C(\rf<10><19> ), .D(
        \rf<11><19> ), .S0(n783), .S1(n768), .Y(n704) );
  OAI2BB2X1 U303 ( .B0(n1028), .B1(n1008), .A0N(N514), .A1N(n1009), .Y(
        \rd1<20> ) );
  MX4X1 U304 ( .A(n710), .B(n708), .C(n709), .D(n707), .S0(n760), .S1(n763), 
        .Y(N514) );
  MX4X1 U305 ( .A(\rf<0><20> ), .B(\rf<1><20> ), .C(\rf<2><20> ), .D(
        \rf<3><20> ), .S0(n783), .S1(n768), .Y(n710) );
  MX4X1 U306 ( .A(\rf<8><20> ), .B(\rf<9><20> ), .C(\rf<10><20> ), .D(
        \rf<11><20> ), .S0(n783), .S1(n768), .Y(n708) );
  OAI2BB2X1 U307 ( .B0(n1010), .B1(n1037), .A0N(N556), .A1N(n1012), .Y(
        \rd2<11> ) );
  MX4X1 U308 ( .A(n838), .B(n836), .C(n837), .D(n835), .S0(n923), .S1(n926), 
        .Y(N556) );
  MX4X1 U309 ( .A(\rf<0><11> ), .B(\rf<1><11> ), .C(\rf<2><11> ), .D(
        \rf<3><11> ), .S0(N16), .S1(n935), .Y(n838) );
  MX4X1 U310 ( .A(\rf<8><11> ), .B(\rf<9><11> ), .C(\rf<10><11> ), .D(
        \rf<11><11> ), .S0(n943), .S1(n935), .Y(n836) );
  OAI2BB2X1 U311 ( .B0(n1011), .B1(n1036), .A0N(N555), .A1N(n1012), .Y(
        \rd2<12> ) );
  MX4X1 U312 ( .A(n842), .B(n840), .C(n841), .D(n839), .S0(n923), .S1(n926), 
        .Y(N555) );
  MX4X1 U313 ( .A(\rf<0><12> ), .B(\rf<1><12> ), .C(\rf<2><12> ), .D(
        \rf<3><12> ), .S0(n949), .S1(n930), .Y(n842) );
  MX4X1 U314 ( .A(\rf<8><12> ), .B(\rf<9><12> ), .C(\rf<10><12> ), .D(
        \rf<11><12> ), .S0(n937), .S1(n935), .Y(n840) );
  OAI2BB2X1 U315 ( .B0(n1010), .B1(n1035), .A0N(N554), .A1N(n1012), .Y(
        \rd2<13> ) );
  MX4X1 U316 ( .A(n846), .B(n844), .C(n845), .D(n843), .S0(n923), .S1(n926), 
        .Y(N554) );
  MX4X1 U317 ( .A(\rf<0><13> ), .B(\rf<1><13> ), .C(\rf<2><13> ), .D(
        \rf<3><13> ), .S0(n943), .S1(n933), .Y(n846) );
  MX4X1 U318 ( .A(\rf<8><13> ), .B(\rf<9><13> ), .C(\rf<10><13> ), .D(
        \rf<11><13> ), .S0(n937), .S1(n931), .Y(n844) );
  OAI2BB2X1 U319 ( .B0(n1011), .B1(n1034), .A0N(N553), .A1N(n1012), .Y(
        \rd2<14> ) );
  MX4X1 U320 ( .A(n850), .B(n848), .C(n849), .D(n847), .S0(n923), .S1(n926), 
        .Y(N553) );
  MX4X1 U321 ( .A(\rf<0><14> ), .B(\rf<1><14> ), .C(\rf<2><14> ), .D(
        \rf<3><14> ), .S0(n948), .S1(N17), .Y(n850) );
  MX4X1 U322 ( .A(\rf<8><14> ), .B(\rf<9><14> ), .C(\rf<10><14> ), .D(
        \rf<11><14> ), .S0(n943), .S1(n931), .Y(n848) );
  OAI2BB2X1 U323 ( .B0(n1010), .B1(n1033), .A0N(N552), .A1N(n1012), .Y(
        \rd2<15> ) );
  MX4X1 U324 ( .A(n854), .B(n852), .C(n853), .D(n851), .S0(n923), .S1(n926), 
        .Y(N552) );
  MX4X1 U325 ( .A(\rf<0><15> ), .B(\rf<1><15> ), .C(\rf<2><15> ), .D(
        \rf<3><15> ), .S0(n945), .S1(n931), .Y(n854) );
  MX4X1 U326 ( .A(\rf<8><15> ), .B(\rf<9><15> ), .C(\rf<10><15> ), .D(
        \rf<11><15> ), .S0(n948), .S1(n932), .Y(n852) );
  OAI2BB2X1 U327 ( .B0(n1037), .B1(n1008), .A0N(N523), .A1N(n1009), .Y(
        \rd1<11> ) );
  MX4X1 U328 ( .A(n674), .B(n672), .C(n673), .D(n671), .S0(n759), .S1(n762), 
        .Y(N523) );
  MX4X1 U329 ( .A(\rf<0><11> ), .B(\rf<1><11> ), .C(\rf<2><11> ), .D(
        \rf<3><11> ), .S0(n786), .S1(n771), .Y(n674) );
  MX4X1 U330 ( .A(\rf<8><11> ), .B(\rf<9><11> ), .C(\rf<10><11> ), .D(
        \rf<11><11> ), .S0(n786), .S1(n771), .Y(n672) );
  OAI2BB2X1 U331 ( .B0(n1036), .B1(n1007), .A0N(N522), .A1N(n1009), .Y(
        \rd1<12> ) );
  MX4X1 U332 ( .A(n678), .B(n676), .C(n677), .D(n675), .S0(n759), .S1(n762), 
        .Y(N522) );
  MX4X1 U333 ( .A(\rf<0><12> ), .B(\rf<1><12> ), .C(\rf<2><12> ), .D(
        \rf<3><12> ), .S0(n785), .S1(n770), .Y(n678) );
  MX4X1 U334 ( .A(\rf<8><12> ), .B(\rf<9><12> ), .C(\rf<10><12> ), .D(
        \rf<11><12> ), .S0(n786), .S1(n771), .Y(n676) );
  OAI2BB2X1 U335 ( .B0(n1035), .B1(n1008), .A0N(N521), .A1N(n1009), .Y(
        \rd1<13> ) );
  MX4X1 U336 ( .A(n682), .B(n680), .C(n681), .D(n679), .S0(n759), .S1(n762), 
        .Y(N521) );
  MX4X1 U337 ( .A(\rf<0><13> ), .B(\rf<1><13> ), .C(\rf<2><13> ), .D(
        \rf<3><13> ), .S0(n785), .S1(n770), .Y(n682) );
  MX4X1 U338 ( .A(\rf<8><13> ), .B(\rf<9><13> ), .C(\rf<10><13> ), .D(
        \rf<11><13> ), .S0(n785), .S1(n770), .Y(n680) );
  OAI2BB2X1 U339 ( .B0(n1034), .B1(n1007), .A0N(N520), .A1N(n1009), .Y(
        \rd1<14> ) );
  MX4X1 U340 ( .A(n686), .B(n684), .C(n685), .D(n683), .S0(n759), .S1(n762), 
        .Y(N520) );
  MX4X1 U341 ( .A(\rf<0><14> ), .B(\rf<1><14> ), .C(\rf<2><14> ), .D(
        \rf<3><14> ), .S0(n785), .S1(n770), .Y(n686) );
  MX4X1 U342 ( .A(\rf<8><14> ), .B(\rf<9><14> ), .C(\rf<10><14> ), .D(
        \rf<11><14> ), .S0(n785), .S1(n770), .Y(n684) );
  OAI2BB2X1 U343 ( .B0(n1033), .B1(n1008), .A0N(N519), .A1N(n1009), .Y(
        \rd1<15> ) );
  MX4X1 U344 ( .A(n690), .B(n688), .C(n689), .D(n687), .S0(n759), .S1(n762), 
        .Y(N519) );
  MX4X1 U345 ( .A(\rf<0><15> ), .B(\rf<1><15> ), .C(\rf<2><15> ), .D(
        \rf<3><15> ), .S0(n785), .S1(n770), .Y(n690) );
  MX4X1 U346 ( .A(\rf<8><15> ), .B(\rf<9><15> ), .C(\rf<10><15> ), .D(
        \rf<11><15> ), .S0(n785), .S1(n770), .Y(n688) );
  OAI2BB2X1 U347 ( .B0(n1010), .B1(n1042), .A0N(N561), .A1N(n1011), .Y(
        \rd2<6> ) );
  MX4X1 U348 ( .A(n818), .B(n816), .C(n817), .D(n815), .S0(n923), .S1(n926), 
        .Y(N561) );
  MX4X1 U349 ( .A(\rf<0><6> ), .B(\rf<1><6> ), .C(\rf<2><6> ), .D(\rf<3><6> ), 
        .S0(n947), .S1(n929), .Y(n818) );
  MX4X1 U350 ( .A(\rf<8><6> ), .B(\rf<9><6> ), .C(\rf<10><6> ), .D(\rf<11><6> ), .S0(n948), .S1(n934), .Y(n816) );
  OAI2BB2X1 U351 ( .B0(n1010), .B1(n1041), .A0N(N560), .A1N(n1012), .Y(
        \rd2<7> ) );
  MX4X1 U352 ( .A(n822), .B(n820), .C(n821), .D(n819), .S0(n923), .S1(n927), 
        .Y(N560) );
  MX4X1 U353 ( .A(\rf<0><7> ), .B(\rf<1><7> ), .C(\rf<2><7> ), .D(\rf<3><7> ), 
        .S0(n946), .S1(n934), .Y(n822) );
  MX4X1 U354 ( .A(\rf<8><7> ), .B(\rf<9><7> ), .C(\rf<10><7> ), .D(\rf<11><7> ), .S0(n945), .S1(n935), .Y(n820) );
  OAI2BB2X1 U355 ( .B0(n1010), .B1(n1040), .A0N(N559), .A1N(n1010), .Y(
        \rd2<8> ) );
  MX4X1 U356 ( .A(n826), .B(n824), .C(n825), .D(n823), .S0(n923), .S1(n926), 
        .Y(N559) );
  MX4X1 U357 ( .A(\rf<0><8> ), .B(\rf<1><8> ), .C(\rf<2><8> ), .D(\rf<3><8> ), 
        .S0(n944), .S1(n932), .Y(n826) );
  MX4X1 U358 ( .A(\rf<8><8> ), .B(\rf<9><8> ), .C(\rf<10><8> ), .D(\rf<11><8> ), .S0(n949), .S1(N17), .Y(n824) );
  OAI2BB2X1 U359 ( .B0(n1011), .B1(n1039), .A0N(N558), .A1N(n1010), .Y(
        \rd2<9> ) );
  MX4X1 U360 ( .A(n830), .B(n828), .C(n829), .D(n827), .S0(n923), .S1(n926), 
        .Y(N558) );
  MX4X1 U361 ( .A(\rf<0><9> ), .B(\rf<1><9> ), .C(\rf<2><9> ), .D(\rf<3><9> ), 
        .S0(n944), .S1(n935), .Y(n830) );
  MX4X1 U362 ( .A(\rf<8><9> ), .B(\rf<9><9> ), .C(\rf<10><9> ), .D(\rf<11><9> ), .S0(n948), .S1(n934), .Y(n828) );
  OAI2BB2X1 U363 ( .B0(n1011), .B1(n1038), .A0N(N557), .A1N(n1012), .Y(
        \rd2<10> ) );
  MX4X1 U364 ( .A(n834), .B(n832), .C(n833), .D(n831), .S0(n923), .S1(n926), 
        .Y(N557) );
  MX4X1 U365 ( .A(\rf<0><10> ), .B(\rf<1><10> ), .C(\rf<2><10> ), .D(
        \rf<3><10> ), .S0(n944), .S1(n935), .Y(n834) );
  MX4X1 U366 ( .A(\rf<8><10> ), .B(\rf<9><10> ), .C(\rf<10><10> ), .D(
        \rf<11><10> ), .S0(n937), .S1(n935), .Y(n832) );
  OAI2BB2X1 U367 ( .B0(n1042), .B1(n1007), .A0N(N528), .A1N(n1009), .Y(
        \rd1<6> ) );
  MX4X1 U368 ( .A(n654), .B(n652), .C(n653), .D(n651), .S0(n759), .S1(N14), 
        .Y(N528) );
  MX4X1 U369 ( .A(\rf<0><6> ), .B(\rf<1><6> ), .C(\rf<2><6> ), .D(\rf<3><6> ), 
        .S0(n787), .S1(n772), .Y(n654) );
  MX4X1 U370 ( .A(\rf<8><6> ), .B(\rf<9><6> ), .C(\rf<10><6> ), .D(\rf<11><6> ), .S0(n783), .S1(n768), .Y(n652) );
  OAI2BB2X1 U371 ( .B0(n1041), .B1(n1007), .A0N(N527), .A1N(n1009), .Y(
        \rd1<7> ) );
  MX4X1 U372 ( .A(n658), .B(n656), .C(n657), .D(n655), .S0(n760), .S1(n763), 
        .Y(N527) );
  MX4X1 U373 ( .A(\rf<0><7> ), .B(\rf<1><7> ), .C(\rf<2><7> ), .D(\rf<3><7> ), 
        .S0(n787), .S1(n768), .Y(n658) );
  MX4X1 U374 ( .A(\rf<8><7> ), .B(\rf<9><7> ), .C(\rf<10><7> ), .D(\rf<11><7> ), .S0(n787), .S1(n772), .Y(n656) );
  OAI2BB2X1 U375 ( .B0(n1040), .B1(n1007), .A0N(N526), .A1N(n1009), .Y(
        \rd1<8> ) );
  MX4X1 U376 ( .A(n662), .B(n660), .C(n661), .D(n659), .S0(n759), .S1(n762), 
        .Y(N526) );
  MX4X1 U377 ( .A(\rf<0><8> ), .B(\rf<1><8> ), .C(\rf<2><8> ), .D(\rf<3><8> ), 
        .S0(n787), .S1(n767), .Y(n662) );
  MX4X1 U378 ( .A(\rf<8><8> ), .B(\rf<9><8> ), .C(\rf<10><8> ), .D(\rf<11><8> ), .S0(n787), .S1(n772), .Y(n660) );
  OAI2BB2X1 U379 ( .B0(n1039), .B1(n1008), .A0N(N525), .A1N(n1007), .Y(
        \rd1<9> ) );
  MX4X1 U380 ( .A(n666), .B(n664), .C(n665), .D(n663), .S0(n759), .S1(n762), 
        .Y(N525) );
  MX4X1 U381 ( .A(\rf<0><9> ), .B(\rf<1><9> ), .C(\rf<2><9> ), .D(\rf<3><9> ), 
        .S0(n786), .S1(n771), .Y(n666) );
  MX4X1 U382 ( .A(\rf<8><9> ), .B(\rf<9><9> ), .C(\rf<10><9> ), .D(\rf<11><9> ), .S0(n787), .S1(n772), .Y(n664) );
  OAI2BB2X1 U383 ( .B0(n1038), .B1(n1007), .A0N(N524), .A1N(n1009), .Y(
        \rd1<10> ) );
  MX4X1 U384 ( .A(n670), .B(n668), .C(n669), .D(n667), .S0(n759), .S1(n762), 
        .Y(N524) );
  MX4X1 U385 ( .A(\rf<0><10> ), .B(\rf<1><10> ), .C(\rf<2><10> ), .D(
        \rf<3><10> ), .S0(n786), .S1(n771), .Y(n670) );
  MX4X1 U386 ( .A(\rf<8><10> ), .B(\rf<9><10> ), .C(\rf<10><10> ), .D(
        \rf<11><10> ), .S0(n786), .S1(n771), .Y(n668) );
  OAI2BB2X1 U387 ( .B0(n1011), .B1(n1047), .A0N(N566), .A1N(n1011), .Y(
        \rd2<1> ) );
  MX4X1 U388 ( .A(n798), .B(n796), .C(n797), .D(n795), .S0(n924), .S1(n926), 
        .Y(N566) );
  MX4X1 U389 ( .A(\rf<0><1> ), .B(\rf<1><1> ), .C(\rf<2><1> ), .D(\rf<3><1> ), 
        .S0(n947), .S1(n933), .Y(n798) );
  MX4X1 U390 ( .A(\rf<8><1> ), .B(\rf<9><1> ), .C(\rf<10><1> ), .D(\rf<11><1> ), .S0(n946), .S1(n932), .Y(n796) );
  OAI2BB2X1 U391 ( .B0(n1010), .B1(n1046), .A0N(N565), .A1N(n1012), .Y(
        \rd2<2> ) );
  MX4X1 U392 ( .A(n802), .B(n800), .C(n801), .D(n799), .S0(n923), .S1(n926), 
        .Y(N565) );
  MX4X1 U393 ( .A(\rf<0><2> ), .B(\rf<1><2> ), .C(\rf<2><2> ), .D(\rf<3><2> ), 
        .S0(n948), .S1(n934), .Y(n802) );
  MX4X1 U394 ( .A(\rf<8><2> ), .B(\rf<9><2> ), .C(\rf<10><2> ), .D(\rf<11><2> ), .S0(n947), .S1(n933), .Y(n800) );
  OAI2BB2X1 U395 ( .B0(n1010), .B1(n1045), .A0N(N564), .A1N(n1010), .Y(
        \rd2<3> ) );
  MX4X1 U396 ( .A(n806), .B(n804), .C(n805), .D(n803), .S0(n923), .S1(n927), 
        .Y(N564) );
  MX4X1 U397 ( .A(\rf<0><3> ), .B(\rf<1><3> ), .C(\rf<2><3> ), .D(\rf<3><3> ), 
        .S0(n949), .S1(n933), .Y(n806) );
  MX4X1 U398 ( .A(\rf<8><3> ), .B(\rf<9><3> ), .C(\rf<10><3> ), .D(\rf<11><3> ), .S0(n949), .S1(n931), .Y(n804) );
  OAI2BB2X1 U399 ( .B0(n1010), .B1(n1044), .A0N(N563), .A1N(n1011), .Y(
        \rd2<4> ) );
  MX4X1 U400 ( .A(n810), .B(n808), .C(n809), .D(n807), .S0(n924), .S1(n926), 
        .Y(N563) );
  MX4X1 U401 ( .A(\rf<0><4> ), .B(\rf<1><4> ), .C(\rf<2><4> ), .D(\rf<3><4> ), 
        .S0(N16), .S1(n935), .Y(n810) );
  MX4X1 U402 ( .A(\rf<8><4> ), .B(\rf<9><4> ), .C(\rf<10><4> ), .D(\rf<11><4> ), .S0(n946), .S1(n930), .Y(n808) );
  OAI2BB2X1 U403 ( .B0(n1010), .B1(n1043), .A0N(N562), .A1N(n1012), .Y(
        \rd2<5> ) );
  MX4X1 U404 ( .A(n814), .B(n812), .C(n813), .D(n811), .S0(n924), .S1(n927), 
        .Y(N562) );
  MX4X1 U405 ( .A(\rf<0><5> ), .B(\rf<1><5> ), .C(\rf<2><5> ), .D(\rf<3><5> ), 
        .S0(n949), .S1(n935), .Y(n814) );
  MX4X1 U406 ( .A(\rf<8><5> ), .B(\rf<9><5> ), .C(\rf<10><5> ), .D(\rf<11><5> ), .S0(N16), .S1(n935), .Y(n812) );
  OAI2BB2X1 U407 ( .B0(n1047), .B1(n1008), .A0N(N533), .A1N(n1007), .Y(
        \rd1<1> ) );
  MX4X1 U408 ( .A(n634), .B(n632), .C(n633), .D(n631), .S0(N15), .S1(N14), .Y(
        N533) );
  MX4X1 U409 ( .A(\rf<0><1> ), .B(\rf<1><1> ), .C(\rf<2><1> ), .D(\rf<3><1> ), 
        .S0(n782), .S1(n768), .Y(n634) );
  MX4X1 U410 ( .A(\rf<8><1> ), .B(\rf<9><1> ), .C(\rf<10><1> ), .D(\rf<11><1> ), .S0(n781), .S1(n767), .Y(n632) );
  OAI2BB2X1 U411 ( .B0(n1046), .B1(n1007), .A0N(N532), .A1N(n1009), .Y(
        \rd1<2> ) );
  MX4X1 U412 ( .A(n638), .B(n636), .C(n637), .D(n635), .S0(n759), .S1(n762), 
        .Y(N532) );
  MX4X1 U413 ( .A(\rf<0><2> ), .B(\rf<1><2> ), .C(\rf<2><2> ), .D(\rf<3><2> ), 
        .S0(n783), .S1(n768), .Y(n638) );
  MX4X1 U414 ( .A(\rf<8><2> ), .B(\rf<9><2> ), .C(\rf<10><2> ), .D(\rf<11><2> ), .S0(n782), .S1(N13), .Y(n636) );
  OAI2BB2X1 U415 ( .B0(n1045), .B1(n1007), .A0N(N531), .A1N(n1008), .Y(
        \rd1<3> ) );
  MX4X1 U416 ( .A(n642), .B(n640), .C(n641), .D(n639), .S0(N15), .S1(n762), 
        .Y(N531) );
  MX4X1 U417 ( .A(\rf<0><3> ), .B(\rf<1><3> ), .C(\rf<2><3> ), .D(\rf<3><3> ), 
        .S0(n784), .S1(n769), .Y(n642) );
  MX4X1 U418 ( .A(\rf<8><3> ), .B(\rf<9><3> ), .C(\rf<10><3> ), .D(\rf<11><3> ), .S0(n784), .S1(n769), .Y(n640) );
  OAI2BB2X1 U419 ( .B0(n1044), .B1(n1007), .A0N(N530), .A1N(n1007), .Y(
        \rd1<4> ) );
  MX4X1 U420 ( .A(n646), .B(n644), .C(n645), .D(n643), .S0(N15), .S1(N14), .Y(
        N530) );
  MX4X1 U421 ( .A(\rf<0><4> ), .B(\rf<1><4> ), .C(\rf<2><4> ), .D(\rf<3><4> ), 
        .S0(n786), .S1(n771), .Y(n646) );
  MX4X1 U422 ( .A(\rf<8><4> ), .B(\rf<9><4> ), .C(\rf<10><4> ), .D(\rf<11><4> ), .S0(n785), .S1(n770), .Y(n644) );
  OAI2BB2X1 U423 ( .B0(n1043), .B1(n1007), .A0N(N529), .A1N(n1008), .Y(
        \rd1<5> ) );
  MX4X1 U424 ( .A(n650), .B(n648), .C(n649), .D(n647), .S0(N15), .S1(N14), .Y(
        N529) );
  MX4X1 U425 ( .A(\rf<0><5> ), .B(\rf<1><5> ), .C(\rf<2><5> ), .D(\rf<3><5> ), 
        .S0(n787), .S1(n765), .Y(n650) );
  MX4X1 U426 ( .A(\rf<8><5> ), .B(\rf<9><5> ), .C(\rf<10><5> ), .D(\rf<11><5> ), .S0(n786), .S1(n771), .Y(n648) );
  OAI2BB2X1 U427 ( .B0(n1010), .B1(n1048), .A0N(N567), .A1N(n1012), .Y(
        \rd2<0> ) );
  MX4X1 U428 ( .A(n794), .B(n792), .C(n793), .D(n791), .S0(n923), .S1(n927), 
        .Y(N567) );
  MX4X1 U429 ( .A(\rf<0><0> ), .B(\rf<1><0> ), .C(\rf<2><0> ), .D(\rf<3><0> ), 
        .S0(n946), .S1(n932), .Y(n794) );
  MX4X1 U430 ( .A(\rf<8><0> ), .B(\rf<9><0> ), .C(\rf<10><0> ), .D(\rf<11><0> ), .S0(n945), .S1(n931), .Y(n792) );
  OAI2BB2X1 U431 ( .B0(n1048), .B1(n1008), .A0N(N534), .A1N(n1009), .Y(
        \rd1<0> ) );
  MX4X1 U432 ( .A(n630), .B(n628), .C(n629), .D(n627), .S0(n760), .S1(n763), 
        .Y(N534) );
  MX4X1 U433 ( .A(\rf<0><0> ), .B(\rf<1><0> ), .C(\rf<2><0> ), .D(\rf<3><0> ), 
        .S0(n781), .S1(n765), .Y(n630) );
  MX4X1 U434 ( .A(\rf<8><0> ), .B(\rf<9><0> ), .C(\rf<10><0> ), .D(\rf<11><0> ), .S0(n784), .S1(n767), .Y(n628) );
  MX4X1 U435 ( .A(\rf<4><0> ), .B(\rf<5><0> ), .C(\rf<6><0> ), .D(\rf<7><0> ), 
        .S0(n783), .S1(n767), .Y(n629) );
  MX4X1 U436 ( .A(\rf<4><1> ), .B(\rf<5><1> ), .C(\rf<6><1> ), .D(\rf<7><1> ), 
        .S0(n782), .S1(n765), .Y(n633) );
  MX4X1 U437 ( .A(\rf<4><2> ), .B(\rf<5><2> ), .C(\rf<6><2> ), .D(\rf<7><2> ), 
        .S0(n783), .S1(n768), .Y(n637) );
  MX4X1 U438 ( .A(\rf<4><3> ), .B(\rf<5><3> ), .C(\rf<6><3> ), .D(\rf<7><3> ), 
        .S0(n784), .S1(n769), .Y(n641) );
  MX4X1 U439 ( .A(\rf<4><4> ), .B(\rf<5><4> ), .C(\rf<6><4> ), .D(\rf<7><4> ), 
        .S0(n785), .S1(n770), .Y(n645) );
  MX4X1 U440 ( .A(\rf<4><5> ), .B(\rf<5><5> ), .C(\rf<6><5> ), .D(\rf<7><5> ), 
        .S0(n787), .S1(n771), .Y(n649) );
  MX4X1 U441 ( .A(\rf<4><6> ), .B(\rf<5><6> ), .C(\rf<6><6> ), .D(\rf<7><6> ), 
        .S0(n787), .S1(n770), .Y(n653) );
  MX4X1 U442 ( .A(\rf<4><7> ), .B(\rf<5><7> ), .C(\rf<6><7> ), .D(\rf<7><7> ), 
        .S0(n787), .S1(n769), .Y(n657) );
  MX4X1 U443 ( .A(\rf<4><8> ), .B(\rf<5><8> ), .C(\rf<6><8> ), .D(\rf<7><8> ), 
        .S0(n787), .S1(n768), .Y(n661) );
  MX4X1 U444 ( .A(\rf<4><9> ), .B(\rf<5><9> ), .C(\rf<6><9> ), .D(\rf<7><9> ), 
        .S0(n786), .S1(n771), .Y(n665) );
  MX4X1 U445 ( .A(\rf<4><10> ), .B(\rf<5><10> ), .C(\rf<6><10> ), .D(
        \rf<7><10> ), .S0(n786), .S1(n771), .Y(n669) );
  MX4X1 U446 ( .A(\rf<4><11> ), .B(\rf<5><11> ), .C(\rf<6><11> ), .D(
        \rf<7><11> ), .S0(n786), .S1(n771), .Y(n673) );
  MX4X1 U447 ( .A(\rf<4><12> ), .B(\rf<5><12> ), .C(\rf<6><12> ), .D(
        \rf<7><12> ), .S0(n786), .S1(n771), .Y(n677) );
  MX4X1 U448 ( .A(\rf<4><13> ), .B(\rf<5><13> ), .C(\rf<6><13> ), .D(
        \rf<7><13> ), .S0(n785), .S1(n770), .Y(n681) );
  MX4X1 U449 ( .A(\rf<4><14> ), .B(\rf<5><14> ), .C(\rf<6><14> ), .D(
        \rf<7><14> ), .S0(n785), .S1(n770), .Y(n685) );
  MX4X1 U450 ( .A(\rf<4><15> ), .B(\rf<5><15> ), .C(\rf<6><15> ), .D(
        \rf<7><15> ), .S0(n785), .S1(n770), .Y(n689) );
  MX4X1 U451 ( .A(\rf<4><16> ), .B(\rf<5><16> ), .C(\rf<6><16> ), .D(
        \rf<7><16> ), .S0(n784), .S1(n769), .Y(n693) );
  MX4X1 U452 ( .A(\rf<4><17> ), .B(\rf<5><17> ), .C(\rf<6><17> ), .D(
        \rf<7><17> ), .S0(n784), .S1(n769), .Y(n697) );
  MX4X1 U453 ( .A(\rf<4><18> ), .B(\rf<5><18> ), .C(\rf<6><18> ), .D(
        \rf<7><18> ), .S0(n784), .S1(n769), .Y(n701) );
  MX4X1 U454 ( .A(\rf<4><19> ), .B(\rf<5><19> ), .C(\rf<6><19> ), .D(
        \rf<7><19> ), .S0(n783), .S1(n768), .Y(n705) );
  MX4X1 U455 ( .A(\rf<4><20> ), .B(\rf<5><20> ), .C(\rf<6><20> ), .D(
        \rf<7><20> ), .S0(n783), .S1(n768), .Y(n709) );
  MX4X1 U456 ( .A(\rf<4><21> ), .B(\rf<5><21> ), .C(\rf<6><21> ), .D(
        \rf<7><21> ), .S0(n783), .S1(n768), .Y(n713) );
  MX4X1 U457 ( .A(\rf<4><22> ), .B(\rf<5><22> ), .C(\rf<6><22> ), .D(
        \rf<7><22> ), .S0(n782), .S1(N13), .Y(n717) );
  MX4X1 U458 ( .A(\rf<4><23> ), .B(\rf<5><23> ), .C(\rf<6><23> ), .D(
        \rf<7><23> ), .S0(n782), .S1(N13), .Y(n721) );
  MX4X1 U459 ( .A(\rf<4><24> ), .B(\rf<5><24> ), .C(\rf<6><24> ), .D(
        \rf<7><24> ), .S0(n782), .S1(N13), .Y(n725) );
  MX4X1 U460 ( .A(\rf<4><25> ), .B(\rf<5><25> ), .C(\rf<6><25> ), .D(
        \rf<7><25> ), .S0(n781), .S1(n766), .Y(n729) );
  MX4X1 U461 ( .A(\rf<4><26> ), .B(\rf<5><26> ), .C(\rf<6><26> ), .D(
        \rf<7><26> ), .S0(n781), .S1(n765), .Y(n733) );
  MX4X1 U462 ( .A(\rf<4><27> ), .B(\rf<5><27> ), .C(\rf<6><27> ), .D(
        \rf<7><27> ), .S0(n781), .S1(n767), .Y(n737) );
  MX4X1 U463 ( .A(\rf<4><28> ), .B(\rf<5><28> ), .C(\rf<6><28> ), .D(
        \rf<7><28> ), .S0(n787), .S1(n767), .Y(n741) );
  MX4X1 U464 ( .A(\rf<4><29> ), .B(\rf<5><29> ), .C(\rf<6><29> ), .D(
        \rf<7><29> ), .S0(n787), .S1(n767), .Y(n747) );
  MX4X1 U465 ( .A(\rf<4><30> ), .B(\rf<5><30> ), .C(\rf<6><30> ), .D(
        \rf<7><30> ), .S0(n783), .S1(n767), .Y(n753) );
  MX4X1 U466 ( .A(\rf<4><31> ), .B(\rf<5><31> ), .C(\rf<6><31> ), .D(
        \rf<7><31> ), .S0(n784), .S1(n767), .Y(n757) );
  MX4X1 U467 ( .A(\rf<4><0> ), .B(\rf<5><0> ), .C(\rf<6><0> ), .D(\rf<7><0> ), 
        .S0(n945), .S1(n931), .Y(n793) );
  MX4X1 U468 ( .A(\rf<4><1> ), .B(\rf<5><1> ), .C(\rf<6><1> ), .D(\rf<7><1> ), 
        .S0(n947), .S1(n933), .Y(n797) );
  MX4X1 U469 ( .A(\rf<4><2> ), .B(\rf<5><2> ), .C(\rf<6><2> ), .D(\rf<7><2> ), 
        .S0(n948), .S1(n934), .Y(n801) );
  MX4X1 U470 ( .A(\rf<4><3> ), .B(\rf<5><3> ), .C(\rf<6><3> ), .D(\rf<7><3> ), 
        .S0(n949), .S1(n934), .Y(n805) );
  MX4X1 U471 ( .A(\rf<4><4> ), .B(\rf<5><4> ), .C(\rf<6><4> ), .D(\rf<7><4> ), 
        .S0(n945), .S1(n930), .Y(n809) );
  MX4X1 U472 ( .A(\rf<4><5> ), .B(\rf<5><5> ), .C(\rf<6><5> ), .D(\rf<7><5> ), 
        .S0(n949), .S1(N17), .Y(n813) );
  MX4X1 U473 ( .A(\rf<4><6> ), .B(\rf<5><6> ), .C(\rf<6><6> ), .D(\rf<7><6> ), 
        .S0(n945), .S1(n932), .Y(n817) );
  MX4X1 U474 ( .A(\rf<4><7> ), .B(\rf<5><7> ), .C(\rf<6><7> ), .D(\rf<7><7> ), 
        .S0(n949), .S1(n933), .Y(n821) );
  MX4X1 U475 ( .A(\rf<4><8> ), .B(\rf<5><8> ), .C(\rf<6><8> ), .D(\rf<7><8> ), 
        .S0(n948), .S1(n931), .Y(n825) );
  MX4X1 U476 ( .A(\rf<4><9> ), .B(\rf<5><9> ), .C(\rf<6><9> ), .D(\rf<7><9> ), 
        .S0(n947), .S1(n935), .Y(n829) );
  MX4X1 U477 ( .A(\rf<4><10> ), .B(\rf<5><10> ), .C(\rf<6><10> ), .D(
        \rf<7><10> ), .S0(n946), .S1(n935), .Y(n833) );
  MX4X1 U478 ( .A(\rf<4><11> ), .B(\rf<5><11> ), .C(\rf<6><11> ), .D(
        \rf<7><11> ), .S0(n943), .S1(n935), .Y(n837) );
  MX4X1 U479 ( .A(\rf<4><12> ), .B(\rf<5><12> ), .C(\rf<6><12> ), .D(
        \rf<7><12> ), .S0(n946), .S1(n935), .Y(n841) );
  MX4X1 U480 ( .A(\rf<4><13> ), .B(\rf<5><13> ), .C(\rf<6><13> ), .D(
        \rf<7><13> ), .S0(n947), .S1(n935), .Y(n845) );
  MX4X1 U481 ( .A(\rf<4><14> ), .B(\rf<5><14> ), .C(\rf<6><14> ), .D(
        \rf<7><14> ), .S0(n947), .S1(n935), .Y(n849) );
  MX4X1 U482 ( .A(\rf<4><15> ), .B(\rf<5><15> ), .C(\rf<6><15> ), .D(
        \rf<7><15> ), .S0(n947), .S1(n935), .Y(n853) );
  MX4X1 U483 ( .A(\rf<4><16> ), .B(\rf<5><16> ), .C(\rf<6><16> ), .D(
        \rf<7><16> ), .S0(n949), .S1(n934), .Y(n857) );
  MX4X1 U484 ( .A(\rf<4><17> ), .B(\rf<5><17> ), .C(\rf<6><17> ), .D(
        \rf<7><17> ), .S0(n949), .S1(n934), .Y(n861) );
  MX4X1 U485 ( .A(\rf<4><18> ), .B(\rf<5><18> ), .C(\rf<6><18> ), .D(
        \rf<7><18> ), .S0(n949), .S1(n934), .Y(n865) );
  MX4X1 U486 ( .A(\rf<4><19> ), .B(\rf<5><19> ), .C(\rf<6><19> ), .D(
        \rf<7><19> ), .S0(n948), .S1(n934), .Y(n869) );
  MX4X1 U487 ( .A(\rf<4><20> ), .B(\rf<5><20> ), .C(\rf<6><20> ), .D(
        \rf<7><20> ), .S0(n948), .S1(n934), .Y(n873) );
  MX4X1 U488 ( .A(\rf<4><21> ), .B(\rf<5><21> ), .C(\rf<6><21> ), .D(
        \rf<7><21> ), .S0(n948), .S1(n934), .Y(n877) );
  MX4X1 U489 ( .A(\rf<4><22> ), .B(\rf<5><22> ), .C(\rf<6><22> ), .D(
        \rf<7><22> ), .S0(n947), .S1(n933), .Y(n881) );
  MX4X1 U490 ( .A(\rf<4><23> ), .B(\rf<5><23> ), .C(\rf<6><23> ), .D(
        \rf<7><23> ), .S0(n947), .S1(n933), .Y(n885) );
  MX4X1 U491 ( .A(\rf<4><24> ), .B(\rf<5><24> ), .C(\rf<6><24> ), .D(
        \rf<7><24> ), .S0(n947), .S1(n933), .Y(n889) );
  MX4X1 U492 ( .A(\rf<4><25> ), .B(\rf<5><25> ), .C(\rf<6><25> ), .D(
        \rf<7><25> ), .S0(n946), .S1(n932), .Y(n893) );
  MX4X1 U493 ( .A(\rf<4><26> ), .B(\rf<5><26> ), .C(\rf<6><26> ), .D(
        \rf<7><26> ), .S0(n946), .S1(n932), .Y(n897) );
  MX4X1 U494 ( .A(\rf<4><27> ), .B(\rf<5><27> ), .C(\rf<6><27> ), .D(
        \rf<7><27> ), .S0(n946), .S1(n932), .Y(n901) );
  MX4X1 U495 ( .A(\rf<4><28> ), .B(\rf<5><28> ), .C(\rf<6><28> ), .D(
        \rf<7><28> ), .S0(n945), .S1(n931), .Y(n905) );
  MX4X1 U496 ( .A(\rf<4><29> ), .B(\rf<5><29> ), .C(\rf<6><29> ), .D(
        \rf<7><29> ), .S0(n945), .S1(n931), .Y(n911) );
  MX4X1 U497 ( .A(\rf<4><30> ), .B(\rf<5><30> ), .C(\rf<6><30> ), .D(
        \rf<7><30> ), .S0(n945), .S1(n931), .Y(n917) );
  MX4X1 U498 ( .A(\rf<4><31> ), .B(\rf<5><31> ), .C(\rf<6><31> ), .D(
        \rf<7><31> ), .S0(n945), .S1(n931), .Y(n921) );
  MX4X1 U499 ( .A(\rf<8><29> ), .B(\rf<9><29> ), .C(\rf<10><29> ), .D(
        \rf<11><29> ), .S0(n781), .S1(n765), .Y(n746) );
  MX4X1 U500 ( .A(\rf<8><30> ), .B(\rf<9><30> ), .C(\rf<10><30> ), .D(
        \rf<11><30> ), .S0(n787), .S1(n767), .Y(n752) );
  MX4X1 U501 ( .A(\rf<8><29> ), .B(\rf<9><29> ), .C(\rf<10><29> ), .D(
        \rf<11><29> ), .S0(n946), .S1(n932), .Y(n910) );
  MX4X1 U502 ( .A(\rf<8><30> ), .B(\rf<9><30> ), .C(\rf<10><30> ), .D(
        \rf<11><30> ), .S0(n945), .S1(n931), .Y(n916) );
  MX2X1 U503 ( .A(\rf<12><29> ), .B(\rf<13><29> ), .S0(n782), .Y(n743) );
  MX2X1 U504 ( .A(\rf<12><30> ), .B(\rf<13><30> ), .S0(n773), .Y(n749) );
  MX2X1 U505 ( .A(\rf<12><29> ), .B(\rf<13><29> ), .S0(n946), .Y(n907) );
  MX2X1 U506 ( .A(\rf<12><30> ), .B(\rf<13><30> ), .S0(n948), .Y(n913) );
  MX2X1 U507 ( .A(n625), .B(n626), .S0(n766), .Y(n627) );
  AND2X2 U508 ( .A(\rf<14><0> ), .B(n777), .Y(n626) );
  MX2X1 U509 ( .A(\rf<12><0> ), .B(\rf<13><0> ), .S0(n784), .Y(n625) );
  MXI2X1 U510 ( .A(n21), .B(n22), .S0(n766), .Y(n631) );
  MXI2X1 U511 ( .A(\rf<12><1> ), .B(\rf<13><1> ), .S0(n785), .Y(n21) );
  NAND2X1 U512 ( .A(\rf<14><1> ), .B(n778), .Y(n22) );
  MXI2X1 U513 ( .A(n23), .B(n24), .S0(n766), .Y(n635) );
  MXI2X1 U514 ( .A(\rf<12><2> ), .B(\rf<13><2> ), .S0(n786), .Y(n23) );
  NAND2X1 U515 ( .A(\rf<14><2> ), .B(n778), .Y(n24) );
  MXI2X1 U516 ( .A(n25), .B(n26), .S0(n766), .Y(n639) );
  MXI2X1 U517 ( .A(\rf<12><3> ), .B(\rf<13><3> ), .S0(n787), .Y(n25) );
  NAND2X1 U518 ( .A(\rf<14><3> ), .B(n776), .Y(n26) );
  MXI2X1 U519 ( .A(n27), .B(n28), .S0(n766), .Y(n643) );
  MXI2X1 U520 ( .A(\rf<12><4> ), .B(\rf<13><4> ), .S0(n781), .Y(n27) );
  NAND2X1 U521 ( .A(\rf<14><4> ), .B(n776), .Y(n28) );
  MXI2X1 U522 ( .A(n29), .B(n30), .S0(n766), .Y(n647) );
  MXI2X1 U523 ( .A(\rf<12><5> ), .B(\rf<13><5> ), .S0(n782), .Y(n29) );
  NAND2X1 U524 ( .A(\rf<14><5> ), .B(n775), .Y(n30) );
  MXI2X1 U525 ( .A(n31), .B(n32), .S0(n766), .Y(n651) );
  MXI2X1 U526 ( .A(\rf<12><6> ), .B(\rf<13><6> ), .S0(n786), .Y(n31) );
  NAND2X1 U527 ( .A(\rf<14><6> ), .B(n776), .Y(n32) );
  MXI2X1 U528 ( .A(n33), .B(n34), .S0(n766), .Y(n655) );
  MXI2X1 U529 ( .A(\rf<12><7> ), .B(\rf<13><7> ), .S0(n784), .Y(n33) );
  NAND2X1 U530 ( .A(\rf<14><7> ), .B(n780), .Y(n34) );
  MXI2X1 U531 ( .A(n35), .B(n36), .S0(n766), .Y(n659) );
  MXI2X1 U532 ( .A(\rf<12><8> ), .B(\rf<13><8> ), .S0(N12), .Y(n35) );
  NAND2X1 U533 ( .A(\rf<14><8> ), .B(n779), .Y(n36) );
  MXI2X1 U534 ( .A(n37), .B(n38), .S0(n766), .Y(n663) );
  MXI2X1 U535 ( .A(\rf<12><9> ), .B(\rf<13><9> ), .S0(N12), .Y(n37) );
  NAND2X1 U536 ( .A(\rf<14><9> ), .B(n775), .Y(n38) );
  MXI2X1 U537 ( .A(n39), .B(n40), .S0(n766), .Y(n667) );
  MXI2X1 U538 ( .A(\rf<12><10> ), .B(\rf<13><10> ), .S0(N12), .Y(n39) );
  NAND2X1 U539 ( .A(\rf<14><10> ), .B(n776), .Y(n40) );
  MXI2X1 U540 ( .A(n41), .B(n42), .S0(n766), .Y(n671) );
  MXI2X1 U541 ( .A(\rf<12><11> ), .B(\rf<13><11> ), .S0(N12), .Y(n41) );
  NAND2X1 U542 ( .A(\rf<14><11> ), .B(n775), .Y(n42) );
  MXI2X1 U543 ( .A(n43), .B(n44), .S0(n765), .Y(n675) );
  MXI2X1 U544 ( .A(\rf<12><12> ), .B(\rf<13><12> ), .S0(n786), .Y(n43) );
  NAND2X1 U545 ( .A(\rf<14><12> ), .B(n775), .Y(n44) );
  MXI2X1 U546 ( .A(n45), .B(n46), .S0(n765), .Y(n679) );
  MXI2X1 U547 ( .A(\rf<12><13> ), .B(\rf<13><13> ), .S0(n781), .Y(n45) );
  NAND2X1 U548 ( .A(\rf<14><13> ), .B(n776), .Y(n46) );
  MXI2X1 U549 ( .A(n47), .B(n48), .S0(n765), .Y(n683) );
  MXI2X1 U550 ( .A(\rf<12><14> ), .B(\rf<13><14> ), .S0(n781), .Y(n47) );
  NAND2X1 U551 ( .A(\rf<14><14> ), .B(n776), .Y(n48) );
  MXI2X1 U552 ( .A(n49), .B(n50), .S0(n765), .Y(n687) );
  MXI2X1 U553 ( .A(\rf<12><15> ), .B(\rf<13><15> ), .S0(n785), .Y(n49) );
  NAND2X1 U554 ( .A(\rf<14><15> ), .B(n777), .Y(n50) );
  MXI2X1 U555 ( .A(n51), .B(n52), .S0(n765), .Y(n691) );
  MXI2X1 U556 ( .A(\rf<12><16> ), .B(\rf<13><16> ), .S0(n781), .Y(n51) );
  NAND2X1 U557 ( .A(\rf<14><16> ), .B(n777), .Y(n52) );
  MXI2X1 U558 ( .A(n53), .B(n54), .S0(n765), .Y(n695) );
  MXI2X1 U559 ( .A(\rf<12><17> ), .B(\rf<13><17> ), .S0(n782), .Y(n53) );
  NAND2X1 U560 ( .A(\rf<14><17> ), .B(n778), .Y(n54) );
  MXI2X1 U561 ( .A(n55), .B(n56), .S0(n765), .Y(n699) );
  MXI2X1 U562 ( .A(\rf<12><18> ), .B(\rf<13><18> ), .S0(n773), .Y(n55) );
  NAND2X1 U563 ( .A(\rf<14><18> ), .B(n778), .Y(n56) );
  MXI2X1 U564 ( .A(n57), .B(n58), .S0(n765), .Y(n703) );
  MXI2X1 U565 ( .A(\rf<12><19> ), .B(\rf<13><19> ), .S0(n786), .Y(n57) );
  NAND2X1 U566 ( .A(\rf<14><19> ), .B(n775), .Y(n58) );
  MXI2X1 U567 ( .A(n59), .B(n60), .S0(n765), .Y(n707) );
  MXI2X1 U568 ( .A(\rf<12><20> ), .B(\rf<13><20> ), .S0(n785), .Y(n59) );
  NAND2X1 U569 ( .A(\rf<14><20> ), .B(n788), .Y(n60) );
  MXI2X1 U570 ( .A(n61), .B(n62), .S0(n765), .Y(n711) );
  MXI2X1 U571 ( .A(\rf<12><21> ), .B(\rf<13><21> ), .S0(n786), .Y(n61) );
  NAND2X1 U572 ( .A(\rf<14><21> ), .B(n780), .Y(n62) );
  MXI2X1 U573 ( .A(n63), .B(n64), .S0(n765), .Y(n715) );
  MXI2X1 U574 ( .A(\rf<12><22> ), .B(\rf<13><22> ), .S0(n785), .Y(n63) );
  NAND2X1 U575 ( .A(\rf<14><22> ), .B(n777), .Y(n64) );
  MXI2X1 U576 ( .A(n65), .B(n66), .S0(n765), .Y(n719) );
  MXI2X1 U577 ( .A(\rf<12><23> ), .B(\rf<13><23> ), .S0(n774), .Y(n65) );
  NAND2X1 U578 ( .A(\rf<14><23> ), .B(n788), .Y(n66) );
  MXI2X1 U579 ( .A(n67), .B(n68), .S0(n765), .Y(n723) );
  MXI2X1 U580 ( .A(\rf<12><24> ), .B(\rf<13><24> ), .S0(n773), .Y(n67) );
  NAND2X1 U581 ( .A(\rf<14><24> ), .B(n778), .Y(n68) );
  MXI2X1 U582 ( .A(n69), .B(n70), .S0(n766), .Y(n755) );
  MXI2X1 U583 ( .A(\rf<12><31> ), .B(\rf<13><31> ), .S0(n783), .Y(n69) );
  NAND2X1 U584 ( .A(\rf<14><31> ), .B(n779), .Y(n70) );
  MX2X1 U585 ( .A(n789), .B(n790), .S0(n930), .Y(n791) );
  AND2X2 U586 ( .A(\rf<14><0> ), .B(n938), .Y(n790) );
  MX2X1 U587 ( .A(\rf<12><0> ), .B(\rf<13><0> ), .S0(n944), .Y(n789) );
  MXI2X1 U588 ( .A(n71), .B(n72), .S0(n930), .Y(n795) );
  MXI2X1 U589 ( .A(\rf<12><1> ), .B(\rf<13><1> ), .S0(n944), .Y(n71) );
  NAND2X1 U590 ( .A(\rf<14><1> ), .B(n938), .Y(n72) );
  MXI2X1 U591 ( .A(n73), .B(n74), .S0(n930), .Y(n799) );
  MXI2X1 U592 ( .A(\rf<12><2> ), .B(\rf<13><2> ), .S0(n944), .Y(n73) );
  NAND2X1 U593 ( .A(\rf<14><2> ), .B(n938), .Y(n74) );
  MXI2X1 U594 ( .A(n75), .B(n76), .S0(n930), .Y(n803) );
  MXI2X1 U595 ( .A(\rf<12><3> ), .B(\rf<13><3> ), .S0(n944), .Y(n75) );
  NAND2X1 U596 ( .A(\rf<14><3> ), .B(n941), .Y(n76) );
  MXI2X1 U597 ( .A(n77), .B(n78), .S0(n930), .Y(n807) );
  MXI2X1 U598 ( .A(\rf<12><4> ), .B(\rf<13><4> ), .S0(n944), .Y(n77) );
  NAND2X1 U599 ( .A(\rf<14><4> ), .B(n942), .Y(n78) );
  MXI2X1 U600 ( .A(n79), .B(n80), .S0(n930), .Y(n811) );
  MXI2X1 U601 ( .A(\rf<12><5> ), .B(\rf<13><5> ), .S0(n944), .Y(n79) );
  NAND2X1 U602 ( .A(\rf<14><5> ), .B(n939), .Y(n80) );
  MXI2X1 U603 ( .A(n81), .B(n82), .S0(n930), .Y(n815) );
  MXI2X1 U604 ( .A(\rf<12><6> ), .B(\rf<13><6> ), .S0(n944), .Y(n81) );
  NAND2X1 U605 ( .A(\rf<14><6> ), .B(n939), .Y(n82) );
  MXI2X1 U606 ( .A(n83), .B(n84), .S0(n930), .Y(n819) );
  MXI2X1 U607 ( .A(\rf<12><7> ), .B(\rf<13><7> ), .S0(n944), .Y(n83) );
  NAND2X1 U608 ( .A(\rf<14><7> ), .B(n938), .Y(n84) );
  MXI2X1 U609 ( .A(n85), .B(n86), .S0(n930), .Y(n823) );
  MXI2X1 U610 ( .A(\rf<12><8> ), .B(\rf<13><8> ), .S0(n944), .Y(n85) );
  NAND2X1 U611 ( .A(\rf<14><8> ), .B(n939), .Y(n86) );
  MXI2X1 U612 ( .A(n87), .B(n88), .S0(n930), .Y(n827) );
  MXI2X1 U613 ( .A(\rf<12><9> ), .B(\rf<13><9> ), .S0(n944), .Y(n87) );
  NAND2X1 U614 ( .A(\rf<14><9> ), .B(n939), .Y(n88) );
  MXI2X1 U615 ( .A(n89), .B(n90), .S0(n930), .Y(n831) );
  MXI2X1 U616 ( .A(\rf<12><10> ), .B(\rf<13><10> ), .S0(n944), .Y(n89) );
  NAND2X1 U617 ( .A(\rf<14><10> ), .B(n938), .Y(n90) );
  MXI2X1 U618 ( .A(n91), .B(n92), .S0(n930), .Y(n835) );
  MXI2X1 U619 ( .A(\rf<12><11> ), .B(\rf<13><11> ), .S0(n944), .Y(n91) );
  NAND2X1 U620 ( .A(\rf<14><11> ), .B(n939), .Y(n92) );
  MXI2X1 U621 ( .A(n93), .B(n94), .S0(n929), .Y(n839) );
  MXI2X1 U622 ( .A(\rf<12><12> ), .B(\rf<13><12> ), .S0(n944), .Y(n93) );
  NAND2X1 U623 ( .A(\rf<14><12> ), .B(n941), .Y(n94) );
  MXI2X1 U624 ( .A(n95), .B(n96), .S0(n929), .Y(n843) );
  MXI2X1 U625 ( .A(\rf<12><13> ), .B(\rf<13><13> ), .S0(n944), .Y(n95) );
  NAND2X1 U626 ( .A(\rf<14><13> ), .B(n942), .Y(n96) );
  MXI2X1 U627 ( .A(n97), .B(n98), .S0(n929), .Y(n847) );
  MXI2X1 U628 ( .A(\rf<12><14> ), .B(\rf<13><14> ), .S0(n943), .Y(n97) );
  NAND2X1 U629 ( .A(\rf<14><14> ), .B(n940), .Y(n98) );
  MXI2X1 U630 ( .A(n99), .B(n100), .S0(n929), .Y(n851) );
  MXI2X1 U631 ( .A(\rf<12><15> ), .B(\rf<13><15> ), .S0(n943), .Y(n99) );
  NAND2X1 U632 ( .A(\rf<14><15> ), .B(n941), .Y(n100) );
  MXI2X1 U633 ( .A(n101), .B(n102), .S0(n929), .Y(n855) );
  MXI2X1 U634 ( .A(\rf<12><16> ), .B(\rf<13><16> ), .S0(n943), .Y(n101) );
  NAND2X1 U635 ( .A(\rf<14><16> ), .B(n941), .Y(n102) );
  MXI2X1 U636 ( .A(n103), .B(n104), .S0(n929), .Y(n859) );
  MXI2X1 U637 ( .A(\rf<12><17> ), .B(\rf<13><17> ), .S0(n943), .Y(n103) );
  NAND2X1 U638 ( .A(\rf<14><17> ), .B(n940), .Y(n104) );
  MXI2X1 U639 ( .A(n105), .B(n106), .S0(n929), .Y(n863) );
  MXI2X1 U640 ( .A(\rf<12><18> ), .B(\rf<13><18> ), .S0(n943), .Y(n105) );
  NAND2X1 U641 ( .A(\rf<14><18> ), .B(n940), .Y(n106) );
  MXI2X1 U642 ( .A(n107), .B(n108), .S0(n929), .Y(n867) );
  MXI2X1 U643 ( .A(\rf<12><19> ), .B(\rf<13><19> ), .S0(n943), .Y(n107) );
  NAND2X1 U644 ( .A(\rf<14><19> ), .B(n941), .Y(n108) );
  MXI2X1 U645 ( .A(n109), .B(n110), .S0(n929), .Y(n871) );
  MXI2X1 U646 ( .A(\rf<12><20> ), .B(\rf<13><20> ), .S0(n943), .Y(n109) );
  NAND2X1 U647 ( .A(\rf<14><20> ), .B(n941), .Y(n110) );
  MXI2X1 U648 ( .A(n111), .B(n112), .S0(n929), .Y(n875) );
  MXI2X1 U649 ( .A(\rf<12><21> ), .B(\rf<13><21> ), .S0(n943), .Y(n111) );
  NAND2X1 U650 ( .A(\rf<14><21> ), .B(n942), .Y(n112) );
  MXI2X1 U651 ( .A(n113), .B(n114), .S0(n929), .Y(n879) );
  MXI2X1 U652 ( .A(\rf<12><22> ), .B(\rf<13><22> ), .S0(n943), .Y(n113) );
  NAND2X1 U653 ( .A(\rf<14><22> ), .B(n942), .Y(n114) );
  MXI2X1 U654 ( .A(n115), .B(n116), .S0(n929), .Y(n883) );
  MXI2X1 U655 ( .A(\rf<12><23> ), .B(\rf<13><23> ), .S0(n943), .Y(n115) );
  NAND2X1 U656 ( .A(\rf<14><23> ), .B(n942), .Y(n116) );
  MXI2X1 U657 ( .A(n117), .B(n118), .S0(n929), .Y(n887) );
  MXI2X1 U658 ( .A(\rf<12><24> ), .B(\rf<13><24> ), .S0(n943), .Y(n117) );
  NAND2X1 U659 ( .A(\rf<14><24> ), .B(n940), .Y(n118) );
  MXI2X1 U660 ( .A(n119), .B(n120), .S0(n930), .Y(n919) );
  MXI2X1 U661 ( .A(\rf<12><31> ), .B(\rf<13><31> ), .S0(n944), .Y(n119) );
  NAND2X1 U662 ( .A(\rf<14><31> ), .B(n942), .Y(n120) );
  MXI2X1 U663 ( .A(n121), .B(n122), .S0(n765), .Y(n727) );
  MXI2X1 U664 ( .A(\rf<12><25> ), .B(\rf<13><25> ), .S0(n781), .Y(n121) );
  NAND2X1 U665 ( .A(\rf<14><25> ), .B(n780), .Y(n122) );
  MXI2X1 U666 ( .A(n123), .B(n124), .S0(n767), .Y(n731) );
  MXI2X1 U667 ( .A(\rf<12><26> ), .B(\rf<13><26> ), .S0(n782), .Y(n123) );
  NAND2X1 U668 ( .A(\rf<14><26> ), .B(n777), .Y(n124) );
  MXI2X1 U669 ( .A(n125), .B(n126), .S0(n766), .Y(n735) );
  MXI2X1 U670 ( .A(\rf<12><27> ), .B(\rf<13><27> ), .S0(n782), .Y(n125) );
  NAND2X1 U671 ( .A(\rf<14><27> ), .B(n777), .Y(n126) );
  MXI2X1 U672 ( .A(n127), .B(n128), .S0(n766), .Y(n739) );
  MXI2X1 U673 ( .A(\rf<12><28> ), .B(\rf<13><28> ), .S0(n781), .Y(n127) );
  NAND2X1 U674 ( .A(\rf<14><28> ), .B(n780), .Y(n128) );
  MXI2X1 U675 ( .A(n129), .B(n130), .S0(n929), .Y(n891) );
  MXI2X1 U676 ( .A(\rf<12><25> ), .B(\rf<13><25> ), .S0(n943), .Y(n129) );
  NAND2X1 U677 ( .A(\rf<14><25> ), .B(n940), .Y(n130) );
  MXI2X1 U678 ( .A(n131), .B(n132), .S0(n929), .Y(n895) );
  MXI2X1 U679 ( .A(\rf<12><26> ), .B(\rf<13><26> ), .S0(n943), .Y(n131) );
  NAND2X1 U680 ( .A(\rf<14><26> ), .B(n941), .Y(n132) );
  MXI2X1 U681 ( .A(n133), .B(n134), .S0(n929), .Y(n899) );
  MXI2X1 U682 ( .A(\rf<12><27> ), .B(\rf<13><27> ), .S0(n943), .Y(n133) );
  NAND2X1 U683 ( .A(\rf<14><27> ), .B(n940), .Y(n134) );
  MXI2X1 U684 ( .A(n135), .B(n136), .S0(n929), .Y(n903) );
  MXI2X1 U685 ( .A(\rf<12><28> ), .B(\rf<13><28> ), .S0(n943), .Y(n135) );
  NAND2X1 U686 ( .A(\rf<14><28> ), .B(n938), .Y(n136) );
  AND2X2 U687 ( .A(\rf<14><29> ), .B(n778), .Y(n744) );
  AND2X2 U688 ( .A(\rf<14><30> ), .B(n775), .Y(n750) );
  AND2X2 U689 ( .A(\rf<14><29> ), .B(n942), .Y(n908) );
  AND2X2 U690 ( .A(\rf<14><30> ), .B(n939), .Y(n914) );
  NOR2X1 U691 ( .A(n1050), .B(\wa3<1> ), .Y(n537) );
  NOR2X1 U692 ( .A(n1049), .B(\wa3<3> ), .Y(n543) );
  NOR2X1 U693 ( .A(\wa3<2> ), .B(\wa3<3> ), .Y(n534) );
  NOR2X1 U694 ( .A(\wa3<0> ), .B(\wa3<1> ), .Y(n535) );
  AND2X2 U695 ( .A(\wa3<1> ), .B(n1050), .Y(n539) );
  AND2X2 U696 ( .A(\wa3<3> ), .B(n1049), .Y(n548) );
  AND2X2 U697 ( .A(\wa3<1> ), .B(\wa3<0> ), .Y(n541) );
  AND2X2 U698 ( .A(\wa3<3> ), .B(\wa3<2> ), .Y(n553) );
  INVX1 U699 ( .A(\wa3<2> ), .Y(n1049) );
  INVX1 U700 ( .A(\wa3<0> ), .Y(n1050) );
  BUFX3 U701 ( .A(we3), .Y(n976) );
endmodule


module extend ( .Instr({\Instr<23> , \Instr<22> , \Instr<21> , \Instr<20> , 
        \Instr<19> , \Instr<18> , \Instr<17> , \Instr<16> , \Instr<15> , 
        \Instr<14> , \Instr<13> , \Instr<12> , \Instr<11> , \Instr<10> , 
        \Instr<9> , \Instr<8> , \Instr<7> , \Instr<6> , \Instr<5> , \Instr<4> , 
        \Instr<3> , \Instr<2> , \Instr<1> , \Instr<0> }), .ImmSrc({\ImmSrc<1> , 
        \ImmSrc<0> }), .ExtImm({\ExtImm<31> , \ExtImm<30> , \ExtImm<29> , 
        \ExtImm<28> , \ExtImm<27> , \ExtImm<26> , \ExtImm<25> , \ExtImm<24> , 
        \ExtImm<23> , \ExtImm<22> , \ExtImm<21> , \ExtImm<20> , \ExtImm<19> , 
        \ExtImm<18> , \ExtImm<17> , \ExtImm<16> , \ExtImm<15> , \ExtImm<14> , 
        \ExtImm<13> , \ExtImm<12> , \ExtImm<11> , \ExtImm<10> , \ExtImm<9> , 
        \ExtImm<8> , \ExtImm<7> , \ExtImm<6> , \ExtImm<5> , \ExtImm<4> , 
        \ExtImm<3> , \ExtImm<2> , \ExtImm<1> , \ExtImm<0> }) );
  input \Instr<23> , \Instr<22> , \Instr<21> , \Instr<20> , \Instr<19> ,
         \Instr<18> , \Instr<17> , \Instr<16> , \Instr<15> , \Instr<14> ,
         \Instr<13> , \Instr<12> , \Instr<11> , \Instr<10> , \Instr<9> ,
         \Instr<8> , \Instr<7> , \Instr<6> , \Instr<5> , \Instr<4> ,
         \Instr<3> , \Instr<2> , \Instr<1> , \Instr<0> , \ImmSrc<1> ,
         \ImmSrc<0> ;
  output \ExtImm<31> , \ExtImm<30> , \ExtImm<29> , \ExtImm<28> , \ExtImm<27> ,
         \ExtImm<26> , \ExtImm<25> , \ExtImm<24> , \ExtImm<23> , \ExtImm<22> ,
         \ExtImm<21> , \ExtImm<20> , \ExtImm<19> , \ExtImm<18> , \ExtImm<17> ,
         \ExtImm<16> , \ExtImm<15> , \ExtImm<14> , \ExtImm<13> , \ExtImm<12> ,
         \ExtImm<11> , \ExtImm<10> , \ExtImm<9> , \ExtImm<8> , \ExtImm<7> ,
         \ExtImm<6> , \ExtImm<5> , \ExtImm<4> , \ExtImm<3> , \ExtImm<2> ,
         \ExtImm<1> , \ExtImm<0> ;
  wire   n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20,
         n21, n22;

  BUFX12 U2 ( .A(\ImmSrc<1> ), .Y(n8) );
  CLKBUFX4 U3 ( .A(n9), .Y(n7) );
  INVX1 U4 ( .A(\Instr<1> ), .Y(n21) );
  INVX1 U5 ( .A(\Instr<0> ), .Y(n22) );
  INVX1 U6 ( .A(\Instr<2> ), .Y(n20) );
  INVX1 U7 ( .A(\Instr<3> ), .Y(n19) );
  INVX1 U8 ( .A(\Instr<5> ), .Y(n17) );
  INVX1 U9 ( .A(\Instr<4> ), .Y(n18) );
  INVX1 U10 ( .A(\ImmSrc<0> ), .Y(n10) );
  OAI22XL U11 ( .A0(n7), .A1(n22), .B0(n8), .B1(n20), .Y(\ExtImm<2> ) );
  OAI22XL U12 ( .A0(n7), .A1(n20), .B0(n8), .B1(n18), .Y(\ExtImm<4> ) );
  NOR2BXL U13 ( .AN(\Instr<14> ), .B(n7), .Y(\ExtImm<16> ) );
  NOR2BXL U14 ( .AN(\Instr<13> ), .B(n7), .Y(\ExtImm<15> ) );
  NOR2BXL U15 ( .AN(\Instr<12> ), .B(n7), .Y(\ExtImm<14> ) );
  NOR2BXL U16 ( .AN(\Instr<18> ), .B(n7), .Y(\ExtImm<20> ) );
  NOR2BXL U17 ( .AN(\Instr<17> ), .B(n7), .Y(\ExtImm<19> ) );
  NOR2BXL U18 ( .AN(\Instr<16> ), .B(n7), .Y(\ExtImm<18> ) );
  NOR2BXL U19 ( .AN(\Instr<15> ), .B(n7), .Y(\ExtImm<17> ) );
  NOR2BXL U20 ( .AN(\Instr<22> ), .B(n7), .Y(\ExtImm<24> ) );
  NOR2BXL U21 ( .AN(\Instr<21> ), .B(n7), .Y(\ExtImm<23> ) );
  NOR2BXL U22 ( .AN(\Instr<20> ), .B(n7), .Y(\ExtImm<22> ) );
  NOR2BXL U23 ( .AN(\Instr<19> ), .B(n7), .Y(\ExtImm<21> ) );
  INVX1 U24 ( .A(n8), .Y(n9) );
  NOR2X1 U25 ( .A(n8), .B(n22), .Y(\ExtImm<0> ) );
  NOR2X1 U26 ( .A(n8), .B(n21), .Y(\ExtImm<1> ) );
  OAI22X1 U27 ( .A0(n7), .A1(n21), .B0(n8), .B1(n19), .Y(\ExtImm<3> ) );
  OAI22X1 U28 ( .A0(n7), .A1(n19), .B0(n8), .B1(n17), .Y(\ExtImm<5> ) );
  OAI22X1 U29 ( .A0(n7), .A1(n18), .B0(n8), .B1(n16), .Y(\ExtImm<6> ) );
  OAI22X1 U30 ( .A0(n7), .A1(n17), .B0(n8), .B1(n15), .Y(\ExtImm<7> ) );
  OAI22X1 U31 ( .A0(n7), .A1(n16), .B0(n10), .B1(n14), .Y(\ExtImm<8> ) );
  OAI22X1 U32 ( .A0(n7), .A1(n15), .B0(n10), .B1(n13), .Y(\ExtImm<9> ) );
  OAI22X1 U33 ( .A0(n7), .A1(n14), .B0(n10), .B1(n12), .Y(\ExtImm<10> ) );
  OAI22X1 U34 ( .A0(n13), .A1(n7), .B0(n10), .B1(n11), .Y(\ExtImm<11> ) );
  NOR2X1 U35 ( .A(n7), .B(n12), .Y(\ExtImm<12> ) );
  NOR2X1 U36 ( .A(n7), .B(n11), .Y(\ExtImm<13> ) );
  INVX1 U37 ( .A(\Instr<9> ), .Y(n13) );
  INVX1 U38 ( .A(\Instr<6> ), .Y(n16) );
  INVX1 U39 ( .A(\Instr<7> ), .Y(n15) );
  INVX1 U40 ( .A(\Instr<8> ), .Y(n14) );
  INVX1 U41 ( .A(\Instr<10> ), .Y(n12) );
  INVX1 U42 ( .A(\Instr<11> ), .Y(n11) );
  BUFX3 U43 ( .A(\ExtImm<25> ), .Y(\ExtImm<31> ) );
  BUFX3 U44 ( .A(\ExtImm<25> ), .Y(\ExtImm<30> ) );
  BUFX3 U45 ( .A(\ExtImm<25> ), .Y(\ExtImm<29> ) );
  BUFX3 U46 ( .A(\ExtImm<25> ), .Y(\ExtImm<28> ) );
  BUFX3 U47 ( .A(\ExtImm<25> ), .Y(\ExtImm<27> ) );
  BUFX3 U48 ( .A(\ExtImm<25> ), .Y(\ExtImm<26> ) );
  AND2X2 U49 ( .A(\Instr<23> ), .B(n8), .Y(\ExtImm<25> ) );
endmodule


module alu_DW01_sub_0 ( .A({\A<31> , \A<30> , \A<29> , \A<28> , \A<27> , 
        \A<26> , \A<25> , \A<24> , \A<23> , \A<22> , \A<21> , \A<20> , \A<19> , 
        \A<18> , \A<17> , \A<16> , \A<15> , \A<14> , \A<13> , \A<12> , \A<11> , 
        \A<10> , \A<9> , \A<8> , \A<7> , \A<6> , \A<5> , \A<4> , \A<3> , 
        \A<2> , \A<1> , \A<0> }), .B({\B<31> , \B<30> , \B<29> , \B<28> , 
        \B<27> , \B<26> , \B<25> , \B<24> , \B<23> , \B<22> , \B<21> , \B<20> , 
        \B<19> , \B<18> , \B<17> , \B<16> , \B<15> , \B<14> , \B<13> , \B<12> , 
        \B<11> , \B<10> , \B<9> , \B<8> , \B<7> , \B<6> , \B<5> , \B<4> , 
        \B<3> , \B<2> , \B<1> , \B<0> }), CI, .DIFF({\DIFF<31> , \DIFF<30> , 
        \DIFF<29> , \DIFF<28> , \DIFF<27> , \DIFF<26> , \DIFF<25> , \DIFF<24> , 
        \DIFF<23> , \DIFF<22> , \DIFF<21> , \DIFF<20> , \DIFF<19> , \DIFF<18> , 
        \DIFF<17> , \DIFF<16> , \DIFF<15> , \DIFF<14> , \DIFF<13> , \DIFF<12> , 
        \DIFF<11> , \DIFF<10> , \DIFF<9> , \DIFF<8> , \DIFF<7> , \DIFF<6> , 
        \DIFF<5> , \DIFF<4> , \DIFF<3> , \DIFF<2> , \DIFF<1> , \DIFF<0> }), CO
 );
  input \A<31> , \A<30> , \A<29> , \A<28> , \A<27> , \A<26> , \A<25> , \A<24> ,
         \A<23> , \A<22> , \A<21> , \A<20> , \A<19> , \A<18> , \A<17> ,
         \A<16> , \A<15> , \A<14> , \A<13> , \A<12> , \A<11> , \A<10> , \A<9> ,
         \A<8> , \A<7> , \A<6> , \A<5> , \A<4> , \A<3> , \A<2> , \A<1> ,
         \A<0> , \B<31> , \B<30> , \B<29> , \B<28> , \B<27> , \B<26> , \B<25> ,
         \B<24> , \B<23> , \B<22> , \B<21> , \B<20> , \B<19> , \B<18> ,
         \B<17> , \B<16> , \B<15> , \B<14> , \B<13> , \B<12> , \B<11> ,
         \B<10> , \B<9> , \B<8> , \B<7> , \B<6> , \B<5> , \B<4> , \B<3> ,
         \B<2> , \B<1> , \B<0> , CI;
  output \DIFF<31> , \DIFF<30> , \DIFF<29> , \DIFF<28> , \DIFF<27> ,
         \DIFF<26> , \DIFF<25> , \DIFF<24> , \DIFF<23> , \DIFF<22> ,
         \DIFF<21> , \DIFF<20> , \DIFF<19> , \DIFF<18> , \DIFF<17> ,
         \DIFF<16> , \DIFF<15> , \DIFF<14> , \DIFF<13> , \DIFF<12> ,
         \DIFF<11> , \DIFF<10> , \DIFF<9> , \DIFF<8> , \DIFF<7> , \DIFF<6> ,
         \DIFF<5> , \DIFF<4> , \DIFF<3> , \DIFF<2> , \DIFF<1> , \DIFF<0> , CO;
  wire   \carry<31> , \carry<30> , \carry<29> , \carry<28> , \carry<27> ,
         \carry<26> , \carry<25> , \carry<24> , \carry<23> , \carry<22> ,
         \carry<21> , \carry<20> , \carry<19> , \carry<18> , \carry<17> ,
         \carry<16> , \carry<15> , \carry<14> , \carry<13> , \carry<12> ,
         \carry<11> , \carry<10> , \carry<9> , \carry<8> , \carry<7> ,
         \carry<6> , \carry<5> , \carry<4> , \carry<3> , \carry<2> ,
         \carry<1> , n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13,
         n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27,
         n28, n29, n30, n31;

  ADDFX2 U2_13 ( .A(\A<13> ), .B(n18), .CI(\carry<13> ), .CO(\carry<14> ), .S(
        \DIFF<13> ) );
  ADDFX2 U2_12 ( .A(\A<12> ), .B(n19), .CI(\carry<12> ), .CO(\carry<13> ), .S(
        \DIFF<12> ) );
  ADDFX2 U2_11 ( .A(\A<11> ), .B(n20), .CI(\carry<11> ), .CO(\carry<12> ), .S(
        \DIFF<11> ) );
  ADDFX2 U2_10 ( .A(\A<10> ), .B(n21), .CI(\carry<10> ), .CO(\carry<11> ), .S(
        \DIFF<10> ) );
  ADDFX2 U2_9 ( .A(\A<9> ), .B(n22), .CI(\carry<9> ), .CO(\carry<10> ), .S(
        \DIFF<9> ) );
  ADDFX2 U2_8 ( .A(\A<8> ), .B(n23), .CI(\carry<8> ), .CO(\carry<9> ), .S(
        \DIFF<8> ) );
  ADDFX2 U2_7 ( .A(\A<7> ), .B(n24), .CI(\carry<7> ), .CO(\carry<8> ), .S(
        \DIFF<7> ) );
  ADDFX2 U2_5 ( .A(\A<5> ), .B(n26), .CI(\carry<5> ), .CO(\carry<6> ), .S(
        \DIFF<5> ) );
  ADDFX2 U2_4 ( .A(\A<4> ), .B(n27), .CI(\carry<4> ), .CO(\carry<5> ), .S(
        \DIFF<4> ) );
  ADDFX2 U2_2 ( .A(\A<2> ), .B(n29), .CI(\carry<2> ), .CO(\carry<3> ), .S(
        \DIFF<2> ) );
  ADDFHX4 U2_19 ( .A(\A<19> ), .B(n12), .CI(\carry<19> ), .CO(\carry<20> ), 
        .S(\DIFF<19> ) );
  ADDFHX4 U2_20 ( .A(\A<20> ), .B(n11), .CI(\carry<20> ), .CO(\carry<21> ), 
        .S(\DIFF<20> ) );
  ADDFHX4 U2_22 ( .A(\A<22> ), .B(n9), .CI(\carry<22> ), .CO(\carry<23> ), .S(
        \DIFF<22> ) );
  ADDFHX4 U2_23 ( .A(\A<23> ), .B(n8), .CI(\carry<23> ), .CO(\carry<24> ), .S(
        \DIFF<23> ) );
  ADDFHX4 U2_29 ( .A(\A<29> ), .B(n2), .CI(\carry<29> ), .CO(\carry<30> ), .S(
        \DIFF<29> ) );
  ADDFHX4 U2_25 ( .A(\A<25> ), .B(n6), .CI(\carry<25> ), .CO(\carry<26> ), .S(
        \DIFF<25> ) );
  ADDFHX4 U2_26 ( .A(\A<26> ), .B(n5), .CI(\carry<26> ), .CO(\carry<27> ), .S(
        \DIFF<26> ) );
  ADDFHX4 U2_28 ( .A(\A<28> ), .B(n3), .CI(\carry<28> ), .CO(\carry<29> ), .S(
        \DIFF<28> ) );
  ADDFHX2 U2_30 ( .A(\A<30> ), .B(n1), .CI(\carry<30> ), .CO(\carry<31> ), .S(
        \DIFF<30> ) );
  ADDFHX2 U2_27 ( .A(\A<27> ), .B(n4), .CI(\carry<27> ), .CO(\carry<28> ), .S(
        \DIFF<27> ) );
  ADDFHX2 U2_24 ( .A(\A<24> ), .B(n7), .CI(\carry<24> ), .CO(\carry<25> ), .S(
        \DIFF<24> ) );
  ADDFHX2 U2_21 ( .A(\A<21> ), .B(n10), .CI(\carry<21> ), .CO(\carry<22> ), 
        .S(\DIFF<21> ) );
  ADDFHX2 U2_18 ( .A(\A<18> ), .B(n13), .CI(\carry<18> ), .CO(\carry<19> ), 
        .S(\DIFF<18> ) );
  ADDFX2 U2_17 ( .A(\A<17> ), .B(n14), .CI(\carry<17> ), .CO(\carry<18> ), .S(
        \DIFF<17> ) );
  ADDFX2 U2_16 ( .A(\A<16> ), .B(n15), .CI(\carry<16> ), .CO(\carry<17> ), .S(
        \DIFF<16> ) );
  ADDFX2 U2_15 ( .A(\A<15> ), .B(n16), .CI(\carry<15> ), .CO(\carry<16> ), .S(
        \DIFF<15> ) );
  ADDFX2 U2_14 ( .A(\A<14> ), .B(n17), .CI(\carry<14> ), .CO(\carry<15> ), .S(
        \DIFF<14> ) );
  ADDFHX2 U2_1 ( .A(\A<1> ), .B(n30), .CI(\carry<1> ), .CO(\carry<2> ), .S(
        \DIFF<1> ) );
  ADDFHX4 U2_3 ( .A(\A<3> ), .B(n28), .CI(\carry<3> ), .CO(\carry<4> ), .S(
        \DIFF<3> ) );
  ADDFHXL U2_6 ( .A(\A<6> ), .B(n25), .CI(\carry<6> ), .CO(\carry<7> ), .S(
        \DIFF<6> ) );
  INVX1 U1 ( .A(\B<19> ), .Y(n12) );
  INVX1 U2 ( .A(\B<14> ), .Y(n17) );
  INVX1 U3 ( .A(\B<15> ), .Y(n16) );
  INVX1 U4 ( .A(\B<16> ), .Y(n15) );
  INVX1 U5 ( .A(\B<17> ), .Y(n14) );
  INVX1 U6 ( .A(\B<18> ), .Y(n13) );
  OR2X4 U7 ( .A(\A<0> ), .B(n31), .Y(\carry<1> ) );
  INVX1 U8 ( .A(\B<20> ), .Y(n11) );
  INVX1 U9 ( .A(\B<21> ), .Y(n10) );
  INVX1 U10 ( .A(\B<30> ), .Y(n1) );
  INVX1 U11 ( .A(\B<22> ), .Y(n9) );
  INVX1 U12 ( .A(\B<23> ), .Y(n8) );
  INVX1 U13 ( .A(\B<24> ), .Y(n7) );
  INVX1 U14 ( .A(\B<25> ), .Y(n6) );
  INVX1 U15 ( .A(\B<29> ), .Y(n2) );
  INVX1 U16 ( .A(\B<26> ), .Y(n5) );
  XNOR2X1 U17 ( .A(n31), .B(\A<0> ), .Y(\DIFF<0> ) );
  INVXL U18 ( .A(\B<27> ), .Y(n4) );
  INVXL U19 ( .A(\B<28> ), .Y(n3) );
  XNOR3X4 U20 ( .A(\A<31> ), .B(\B<31> ), .C(\carry<31> ), .Y(\DIFF<31> ) );
  INVX1 U21 ( .A(\B<1> ), .Y(n30) );
  INVX1 U22 ( .A(\B<2> ), .Y(n29) );
  INVX1 U23 ( .A(\B<3> ), .Y(n28) );
  INVX1 U24 ( .A(\B<4> ), .Y(n27) );
  INVX1 U25 ( .A(\B<5> ), .Y(n26) );
  INVX1 U26 ( .A(\B<6> ), .Y(n25) );
  INVX1 U27 ( .A(\B<7> ), .Y(n24) );
  INVX1 U28 ( .A(\B<8> ), .Y(n23) );
  INVX1 U29 ( .A(\B<9> ), .Y(n22) );
  INVX1 U30 ( .A(\B<10> ), .Y(n21) );
  INVX1 U31 ( .A(\B<11> ), .Y(n20) );
  INVX1 U32 ( .A(\B<12> ), .Y(n19) );
  INVX1 U33 ( .A(\B<13> ), .Y(n18) );
  INVX1 U34 ( .A(\B<0> ), .Y(n31) );
endmodule


module alu_DW01_add_0 ( .A({\A<32> , \A<31> , \A<30> , \A<29> , \A<28> , 
        \A<27> , \A<26> , \A<25> , \A<24> , \A<23> , \A<22> , \A<21> , \A<20> , 
        \A<19> , \A<18> , \A<17> , \A<16> , \A<15> , \A<14> , \A<13> , \A<12> , 
        \A<11> , \A<10> , \A<9> , \A<8> , \A<7> , \A<6> , \A<5> , \A<4> , 
        \A<3> , \A<2> , \A<1> , \A<0> }), .B({\B<32> , \B<31> , \B<30> , 
        \B<29> , \B<28> , \B<27> , \B<26> , \B<25> , \B<24> , \B<23> , \B<22> , 
        \B<21> , \B<20> , \B<19> , \B<18> , \B<17> , \B<16> , \B<15> , \B<14> , 
        \B<13> , \B<12> , \B<11> , \B<10> , \B<9> , \B<8> , \B<7> , \B<6> , 
        \B<5> , \B<4> , \B<3> , \B<2> , \B<1> , \B<0> }), CI, .SUM({\SUM<32> , 
        \SUM<31> , \SUM<30> , \SUM<29> , \SUM<28> , \SUM<27> , \SUM<26> , 
        \SUM<25> , \SUM<24> , \SUM<23> , \SUM<22> , \SUM<21> , \SUM<20> , 
        \SUM<19> , \SUM<18> , \SUM<17> , \SUM<16> , \SUM<15> , \SUM<14> , 
        \SUM<13> , \SUM<12> , \SUM<11> , \SUM<10> , \SUM<9> , \SUM<8> , 
        \SUM<7> , \SUM<6> , \SUM<5> , \SUM<4> , \SUM<3> , \SUM<2> , \SUM<1> , 
        \SUM<0> }), CO );
  input \A<32> , \A<31> , \A<30> , \A<29> , \A<28> , \A<27> , \A<26> , \A<25> ,
         \A<24> , \A<23> , \A<22> , \A<21> , \A<20> , \A<19> , \A<18> ,
         \A<17> , \A<16> , \A<15> , \A<14> , \A<13> , \A<12> , \A<11> ,
         \A<10> , \A<9> , \A<8> , \A<7> , \A<6> , \A<5> , \A<4> , \A<3> ,
         \A<2> , \A<1> , \A<0> , \B<32> , \B<31> , \B<30> , \B<29> , \B<28> ,
         \B<27> , \B<26> , \B<25> , \B<24> , \B<23> , \B<22> , \B<21> ,
         \B<20> , \B<19> , \B<18> , \B<17> , \B<16> , \B<15> , \B<14> ,
         \B<13> , \B<12> , \B<11> , \B<10> , \B<9> , \B<8> , \B<7> , \B<6> ,
         \B<5> , \B<4> , \B<3> , \B<2> , \B<1> , \B<0> , CI;
  output \SUM<32> , \SUM<31> , \SUM<30> , \SUM<29> , \SUM<28> , \SUM<27> ,
         \SUM<26> , \SUM<25> , \SUM<24> , \SUM<23> , \SUM<22> , \SUM<21> ,
         \SUM<20> , \SUM<19> , \SUM<18> , \SUM<17> , \SUM<16> , \SUM<15> ,
         \SUM<14> , \SUM<13> , \SUM<12> , \SUM<11> , \SUM<10> , \SUM<9> ,
         \SUM<8> , \SUM<7> , \SUM<6> , \SUM<5> , \SUM<4> , \SUM<3> , \SUM<2> ,
         \SUM<1> , \SUM<0> , CO;
  wire   \carry<31> , \carry<30> , \carry<29> , \carry<28> , \carry<27> ,
         \carry<26> , \carry<25> , \carry<24> , \carry<23> , \carry<22> ,
         \carry<21> , \carry<20> , \carry<19> , \carry<18> , \carry<17> ,
         \carry<16> , \carry<15> , \carry<14> , \carry<13> , \carry<12> ,
         \carry<11> , \carry<10> , \carry<9> , \carry<8> , \carry<7> ,
         \carry<6> , \carry<5> , \carry<4> , \carry<3> , \carry<2> ,
         \carry<1> ;

  ADDFX2 U1_13 ( .A(\A<13> ), .B(\B<13> ), .CI(\carry<13> ), .CO(\carry<14> ), 
        .S(\SUM<13> ) );
  ADDFX2 U1_12 ( .A(\A<12> ), .B(\B<12> ), .CI(\carry<12> ), .CO(\carry<13> ), 
        .S(\SUM<12> ) );
  ADDFX2 U1_11 ( .A(\A<11> ), .B(\B<11> ), .CI(\carry<11> ), .CO(\carry<12> ), 
        .S(\SUM<11> ) );
  ADDFX2 U1_10 ( .A(\A<10> ), .B(\B<10> ), .CI(\carry<10> ), .CO(\carry<11> ), 
        .S(\SUM<10> ) );
  ADDFX2 U1_9 ( .A(\A<9> ), .B(\B<9> ), .CI(\carry<9> ), .CO(\carry<10> ), .S(
        \SUM<9> ) );
  ADDFX2 U1_8 ( .A(\A<8> ), .B(\B<8> ), .CI(\carry<8> ), .CO(\carry<9> ), .S(
        \SUM<8> ) );
  ADDFX2 U1_7 ( .A(\A<7> ), .B(\B<7> ), .CI(\carry<7> ), .CO(\carry<8> ), .S(
        \SUM<7> ) );
  ADDFX2 U1_5 ( .A(\A<5> ), .B(\B<5> ), .CI(\carry<5> ), .CO(\carry<6> ), .S(
        \SUM<5> ) );
  ADDFX2 U1_4 ( .A(\A<4> ), .B(\B<4> ), .CI(\carry<4> ), .CO(\carry<5> ), .S(
        \SUM<4> ) );
  ADDFHX4 U1_29 ( .A(\A<29> ), .B(\B<29> ), .CI(\carry<29> ), .CO(\carry<30> ), 
        .S(\SUM<29> ) );
  ADDFX2 U1_28 ( .A(\A<28> ), .B(\B<28> ), .CI(\carry<28> ), .CO(\carry<29> ), 
        .S(\SUM<28> ) );
  ADDFX2 U1_27 ( .A(\A<27> ), .B(\B<27> ), .CI(\carry<27> ), .CO(\carry<28> ), 
        .S(\SUM<27> ) );
  ADDFX2 U1_26 ( .A(\A<26> ), .B(\B<26> ), .CI(\carry<26> ), .CO(\carry<27> ), 
        .S(\SUM<26> ) );
  ADDFX2 U1_25 ( .A(\A<25> ), .B(\B<25> ), .CI(\carry<25> ), .CO(\carry<26> ), 
        .S(\SUM<25> ) );
  ADDFX2 U1_24 ( .A(\A<24> ), .B(\B<24> ), .CI(\carry<24> ), .CO(\carry<25> ), 
        .S(\SUM<24> ) );
  ADDFX2 U1_23 ( .A(\A<23> ), .B(\B<23> ), .CI(\carry<23> ), .CO(\carry<24> ), 
        .S(\SUM<23> ) );
  ADDFX2 U1_22 ( .A(\A<22> ), .B(\B<22> ), .CI(\carry<22> ), .CO(\carry<23> ), 
        .S(\SUM<22> ) );
  ADDFX2 U1_21 ( .A(\A<21> ), .B(\B<21> ), .CI(\carry<21> ), .CO(\carry<22> ), 
        .S(\SUM<21> ) );
  ADDFX2 U1_20 ( .A(\A<20> ), .B(\B<20> ), .CI(\carry<20> ), .CO(\carry<21> ), 
        .S(\SUM<20> ) );
  ADDFX2 U1_19 ( .A(\A<19> ), .B(\B<19> ), .CI(\carry<19> ), .CO(\carry<20> ), 
        .S(\SUM<19> ) );
  ADDFX2 U1_18 ( .A(\A<18> ), .B(\B<18> ), .CI(\carry<18> ), .CO(\carry<19> ), 
        .S(\SUM<18> ) );
  ADDFX2 U1_17 ( .A(\A<17> ), .B(\B<17> ), .CI(\carry<17> ), .CO(\carry<18> ), 
        .S(\SUM<17> ) );
  ADDFX2 U1_16 ( .A(\A<16> ), .B(\B<16> ), .CI(\carry<16> ), .CO(\carry<17> ), 
        .S(\SUM<16> ) );
  ADDFX2 U1_15 ( .A(\A<15> ), .B(\B<15> ), .CI(\carry<15> ), .CO(\carry<16> ), 
        .S(\SUM<15> ) );
  ADDFX2 U1_14 ( .A(\A<14> ), .B(\B<14> ), .CI(\carry<14> ), .CO(\carry<15> ), 
        .S(\SUM<14> ) );
  ADDFX2 U1_1 ( .A(\A<1> ), .B(\B<1> ), .CI(\carry<1> ), .CO(\carry<2> ), .S(
        \SUM<1> ) );
  ADDFX2 U1_31 ( .A(\A<31> ), .B(\B<31> ), .CI(\carry<31> ), .CO(\SUM<32> ), 
        .S(\SUM<31> ) );
  ADDFX2 U1_3 ( .A(\A<3> ), .B(\B<3> ), .CI(\carry<3> ), .CO(\carry<4> ), .S(
        \SUM<3> ) );
  ADDFHX4 U1_30 ( .A(\A<30> ), .B(\B<30> ), .CI(\carry<30> ), .CO(\carry<31> ), 
        .S(\SUM<30> ) );
  ADDFHX4 U1_2 ( .A(\A<2> ), .B(\B<2> ), .CI(\carry<2> ), .CO(\carry<3> ), .S(
        \SUM<2> ) );
  ADDFHX4 U1_6 ( .A(\A<6> ), .B(\B<6> ), .CI(\carry<6> ), .CO(\carry<7> ), .S(
        \SUM<6> ) );
  XOR2X1 U1 ( .A(\B<0> ), .B(\A<0> ), .Y(\SUM<0> ) );
  AND2X2 U2 ( .A(\B<0> ), .B(\A<0> ), .Y(\carry<1> ) );
endmodule


module alu ( .a({\a<31> , \a<30> , \a<29> , \a<28> , \a<27> , \a<26> , \a<25> , 
        \a<24> , \a<23> , \a<22> , \a<21> , \a<20> , \a<19> , \a<18> , \a<17> , 
        \a<16> , \a<15> , \a<14> , \a<13> , \a<12> , \a<11> , \a<10> , \a<9> , 
        \a<8> , \a<7> , \a<6> , \a<5> , \a<4> , \a<3> , \a<2> , \a<1> , \a<0> 
        }), .b({\b<31> , \b<30> , \b<29> , \b<28> , \b<27> , \b<26> , \b<25> , 
        \b<24> , \b<23> , \b<22> , \b<21> , \b<20> , \b<19> , \b<18> , \b<17> , 
        \b<16> , \b<15> , \b<14> , \b<13> , \b<12> , \b<11> , \b<10> , \b<9> , 
        \b<8> , \b<7> , \b<6> , \b<5> , \b<4> , \b<3> , \b<2> , \b<1> , \b<0> 
        }), .ALUControl({\ALUControl<1> , \ALUControl<0> }), .Result({
        \Result<31> , \Result<30> , \Result<29> , \Result<28> , \Result<27> , 
        \Result<26> , \Result<25> , \Result<24> , \Result<23> , \Result<22> , 
        \Result<21> , \Result<20> , \Result<19> , \Result<18> , \Result<17> , 
        \Result<16> , \Result<15> , \Result<14> , \Result<13> , \Result<12> , 
        \Result<11> , \Result<10> , \Result<9> , \Result<8> , \Result<7> , 
        \Result<6> , \Result<5> , \Result<4> , \Result<3> , \Result<2> , 
        \Result<1> , \Result<0> }), .ALUFlags({\ALUFlags<3> , \ALUFlags<2> , 
        \ALUFlags<1> , \ALUFlags<0> }) );
  input \a<31> , \a<30> , \a<29> , \a<28> , \a<27> , \a<26> , \a<25> , \a<24> ,
         \a<23> , \a<22> , \a<21> , \a<20> , \a<19> , \a<18> , \a<17> ,
         \a<16> , \a<15> , \a<14> , \a<13> , \a<12> , \a<11> , \a<10> , \a<9> ,
         \a<8> , \a<7> , \a<6> , \a<5> , \a<4> , \a<3> , \a<2> , \a<1> ,
         \a<0> , \b<31> , \b<30> , \b<29> , \b<28> , \b<27> , \b<26> , \b<25> ,
         \b<24> , \b<23> , \b<22> , \b<21> , \b<20> , \b<19> , \b<18> ,
         \b<17> , \b<16> , \b<15> , \b<14> , \b<13> , \b<12> , \b<11> ,
         \b<10> , \b<9> , \b<8> , \b<7> , \b<6> , \b<5> , \b<4> , \b<3> ,
         \b<2> , \b<1> , \b<0> , \ALUControl<1> , \ALUControl<0> ;
  output \Result<31> , \Result<30> , \Result<29> , \Result<28> , \Result<27> ,
         \Result<26> , \Result<25> , \Result<24> , \Result<23> , \Result<22> ,
         \Result<21> , \Result<20> , \Result<19> , \Result<18> , \Result<17> ,
         \Result<16> , \Result<15> , \Result<14> , \Result<13> , \Result<12> ,
         \Result<11> , \Result<10> , \Result<9> , \Result<8> , \Result<7> ,
         \Result<6> , \Result<5> , \Result<4> , \Result<3> , \Result<2> ,
         \Result<1> , \Result<0> , \ALUFlags<3> , \ALUFlags<2> , \ALUFlags<1> ,
         \ALUFlags<0> ;
  wire   N13, N14, N15, N16, N17, N18, N19, N20, N21, N22, N23, N24, N25, N26,
         N27, N28, N29, N30, N31, N32, N33, N34, N35, N36, N37, N38, N39, N40,
         N41, N42, N43, N44, N45, N46, N47, N48, N49, N50, N51, N52, N53, N54,
         N55, N56, N57, N58, N59, N60, N61, N62, N63, N64, N65, N66, N67, N68,
         N69, N70, N71, N72, N73, N74, N75, N76, N77, N173, n12, n13, n14, n15,
         n16, n17, n18, n20, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n122, n123, n1,
         n2, n3, n4, n5, n9, n10, n11, n19, n121, n124, n125, n126, n127, n128,
         n129, n130, n131, n132, n133, n134, n135, n136, n137;
  assign \ALUFlags<2>  = N173;

  alu_DW01_sub_0 sub_440 ( .A({\a<31> , \a<30> , \a<29> , \a<28> , \a<27> , 
        \a<26> , \a<25> , \a<24> , \a<23> , \a<22> , \a<21> , \a<20> , \a<19> , 
        \a<18> , \a<17> , \a<16> , \a<15> , \a<14> , \a<13> , \a<12> , \a<11> , 
        \a<10> , \a<9> , \a<8> , \a<7> , \a<6> , \a<5> , \a<4> , n4, \a<2> , 
        \a<1> , n2}), .B({\b<31> , \b<30> , \b<29> , \b<28> , \b<27> , \b<26> , 
        \b<25> , \b<24> , \b<23> , \b<22> , \b<21> , \b<20> , \b<19> , \b<18> , 
        \b<17> , \b<16> , \b<15> , \b<14> , \b<13> , \b<12> , \b<11> , \b<10> , 
        \b<9> , \b<8> , \b<7> , \b<6> , \b<5> , \b<4> , n1, \b<2> , n3, \b<0> }), .CI(1'b0), .DIFF({N77, N76, N75, N74, N73, N72, N71, N70, N69, N68, N67, 
        N66, N65, N64, N63, N62, N61, N60, N59, N58, N57, N56, N55, N54, N53, 
        N52, N51, N50, N49, N48, N47, N46}) );
  alu_DW01_add_0 add_439 ( .A({1'b0, \a<31> , \a<30> , \a<29> , \a<28> , 
        \a<27> , \a<26> , \a<25> , \a<24> , \a<23> , \a<22> , \a<21> , \a<20> , 
        \a<19> , \a<18> , \a<17> , \a<16> , \a<15> , \a<14> , \a<13> , \a<12> , 
        \a<11> , \a<10> , \a<9> , \a<8> , \a<7> , \a<6> , \a<5> , \a<4> , n4, 
        \a<2> , \a<1> , n2}), .B({1'b0, \b<31> , \b<30> , \b<29> , \b<28> , 
        \b<27> , \b<26> , \b<25> , \b<24> , \b<23> , \b<22> , \b<21> , \b<20> , 
        \b<19> , \b<18> , \b<17> , \b<16> , \b<15> , \b<14> , \b<13> , \b<12> , 
        \b<11> , \b<10> , \b<9> , \b<8> , \b<7> , \b<6> , \b<5> , \b<4> , n1, 
        \b<2> , n3, \b<0> }), .CI(1'b0), .SUM({N45, N44, N43, N42, N41, N40, 
        N39, N38, N37, N36, N35, N34, N33, N32, N31, N30, N29, N28, N27, N26, 
        N25, N24, N23, N22, N21, N20, N19, N18, N17, N16, N15, N14, N13}) );
  BUFX3 U4 ( .A(\b<3> ), .Y(n1) );
  BUFX20 U5 ( .A(\a<0> ), .Y(n2) );
  BUFX8 U6 ( .A(\b<1> ), .Y(n3) );
  NAND2X4 U7 ( .A(n86), .B(n87), .Y(\Result<28> ) );
  AOI22X4 U8 ( .A0(N74), .A1(n20), .B0(N41), .B1(n124), .Y(n86) );
  NAND2X4 U9 ( .A(n83), .B(n84), .Y(\Result<29> ) );
  AOI22X4 U10 ( .A0(N75), .A1(n20), .B0(N42), .B1(n124), .Y(n83) );
  AOI22X4 U11 ( .A0(N76), .A1(n125), .B0(N43), .B1(n121), .Y(n53) );
  NOR3X4 U12 ( .A(n118), .B(n135), .C(n119), .Y(\ALUFlags<0> ) );
  BUFX3 U13 ( .A(\a<3> ), .Y(n4) );
  NAND2X2 U14 ( .A(n53), .B(n54), .Y(\Result<30> ) );
  OAI221X4 U15 ( .A0(n9), .A1(n10), .B0(n129), .B1(n11), .C0(n123), .Y(
        \Result<31> ) );
  AOI22XL U16 ( .A0(n1), .A1(n52), .B0(n4), .B1(n19), .Y(n51) );
  INVX1 U17 ( .A(\b<31> ), .Y(n10) );
  INVX1 U18 ( .A(\a<31> ), .Y(n11) );
  INVX1 U19 ( .A(n122), .Y(n9) );
  OR2X2 U20 ( .A(\ALUControl<0> ), .B(n135), .Y(n5) );
  AOI22X4 U21 ( .A0(N77), .A1(n20), .B0(N44), .B1(n121), .Y(n123) );
  AOI22XL U22 ( .A0(n3), .A1(n117), .B0(\a<1> ), .B1(n128), .Y(n116) );
  OR4XL U23 ( .A(\Result<16> ), .B(\Result<17> ), .C(\Result<18> ), .D(
        \Result<19> ), .Y(n93) );
  OR4XL U24 ( .A(\Result<1> ), .B(\Result<20> ), .C(\Result<21> ), .D(
        \Result<22> ), .Y(n92) );
  NOR4BX4 U25 ( .AN(n12), .B(n13), .C(n14), .D(n15), .Y(N173) );
  OR4X2 U26 ( .A(\Result<31> ), .B(\Result<0> ), .C(\Result<10> ), .D(
        \Result<11> ), .Y(n15) );
  OR4X2 U27 ( .A(\Result<27> ), .B(\Result<28> ), .C(\Result<29> ), .D(
        \Result<2> ), .Y(n40) );
  OR4X2 U28 ( .A(\Result<23> ), .B(\Result<24> ), .C(\Result<25> ), .D(
        \Result<26> ), .Y(n41) );
  OR4XL U29 ( .A(\Result<6> ), .B(\Result<7> ), .C(\Result<8> ), .D(
        \Result<9> ), .Y(n42) );
  AOI22XL U30 ( .A0(\b<0> ), .A1(n27), .B0(n2), .B1(n128), .Y(n26) );
  CLKINVX3 U31 ( .A(n132), .Y(n128) );
  INVX1 U32 ( .A(n19), .Y(n129) );
  INVX1 U33 ( .A(n134), .Y(n131) );
  INVX1 U34 ( .A(n19), .Y(n133) );
  INVX1 U35 ( .A(n19), .Y(n132) );
  INVX1 U36 ( .A(n134), .Y(n130) );
  CLKINVX3 U37 ( .A(n137), .Y(n136) );
  CLKINVX3 U38 ( .A(n127), .Y(n125) );
  CLKINVX3 U39 ( .A(n5), .Y(n124) );
  CLKINVX3 U40 ( .A(n137), .Y(n135) );
  INVX1 U41 ( .A(\ALUControl<1> ), .Y(n137) );
  CLKINVX3 U42 ( .A(n127), .Y(n126) );
  INVX1 U43 ( .A(n129), .Y(n134) );
  OR4X2 U44 ( .A(n40), .B(n41), .C(n42), .D(n43), .Y(n13) );
  OR4X2 U45 ( .A(\Result<30> ), .B(\Result<3> ), .C(\Result<4> ), .D(
        \Result<5> ), .Y(n43) );
  NOR2X1 U46 ( .A(n92), .B(n93), .Y(n12) );
  CLKINVX3 U47 ( .A(n5), .Y(n121) );
  INVX1 U48 ( .A(n20), .Y(n127) );
  OAI2BB1X1 U49 ( .A0N(\a<31> ), .A1N(n136), .B0(n129), .Y(n122) );
  AOI22X1 U50 ( .A0(\b<30> ), .A1(n55), .B0(\a<30> ), .B1(n19), .Y(n54) );
  OAI2BB1X1 U51 ( .A0N(n135), .A1N(\a<30> ), .B0(n130), .Y(n55) );
  XNOR2X1 U52 ( .A(\a<31> ), .B(\Result<31> ), .Y(n118) );
  NAND2X1 U53 ( .A(n68), .B(n69), .Y(\Result<26> ) );
  AOI22X1 U54 ( .A0(\b<26> ), .A1(n70), .B0(\a<26> ), .B1(n128), .Y(n69) );
  AOI22X1 U55 ( .A0(N72), .A1(n125), .B0(N39), .B1(n124), .Y(n68) );
  OAI2BB1X1 U56 ( .A0N(n136), .A1N(\a<26> ), .B0(n132), .Y(n70) );
  NAND2X1 U57 ( .A(n71), .B(n72), .Y(\Result<25> ) );
  AOI22X1 U58 ( .A0(\b<25> ), .A1(n73), .B0(\a<25> ), .B1(n128), .Y(n72) );
  AOI22X1 U59 ( .A0(N71), .A1(n125), .B0(N38), .B1(n124), .Y(n71) );
  OAI2BB1X1 U60 ( .A0N(n136), .A1N(\a<25> ), .B0(n131), .Y(n73) );
  AOI22X1 U61 ( .A0(\b<29> ), .A1(n85), .B0(\a<29> ), .B1(n128), .Y(n84) );
  OAI2BB1X1 U62 ( .A0N(n136), .A1N(\a<29> ), .B0(n132), .Y(n85) );
  AOI22X1 U63 ( .A0(\b<28> ), .A1(n88), .B0(\a<28> ), .B1(n128), .Y(n87) );
  OAI2BB1X1 U64 ( .A0N(n136), .A1N(\a<28> ), .B0(n132), .Y(n88) );
  NAND2X1 U65 ( .A(n89), .B(n90), .Y(\Result<27> ) );
  AOI22X1 U66 ( .A0(\b<27> ), .A1(n91), .B0(\a<27> ), .B1(n128), .Y(n90) );
  AOI22X1 U67 ( .A0(N73), .A1(n125), .B0(N40), .B1(n124), .Y(n89) );
  OAI2BB1X1 U68 ( .A0N(n136), .A1N(\a<27> ), .B0(n133), .Y(n91) );
  NAND2X1 U69 ( .A(n106), .B(n107), .Y(\Result<22> ) );
  AOI22X1 U70 ( .A0(\b<22> ), .A1(n108), .B0(\a<22> ), .B1(n19), .Y(n107) );
  AOI22X1 U71 ( .A0(N68), .A1(n126), .B0(N35), .B1(n124), .Y(n106) );
  OAI2BB1X1 U72 ( .A0N(n136), .A1N(\a<22> ), .B0(n130), .Y(n108) );
  NAND2X1 U73 ( .A(n109), .B(n110), .Y(\Result<21> ) );
  AOI22X1 U74 ( .A0(\b<21> ), .A1(n111), .B0(\a<21> ), .B1(n134), .Y(n110) );
  AOI22X1 U75 ( .A0(N67), .A1(n125), .B0(N34), .B1(n124), .Y(n109) );
  OAI2BB1X1 U76 ( .A0N(n136), .A1N(\a<21> ), .B0(n130), .Y(n111) );
  NAND2X1 U77 ( .A(n112), .B(n113), .Y(\Result<20> ) );
  AOI22X1 U78 ( .A0(\b<20> ), .A1(n114), .B0(\a<20> ), .B1(n128), .Y(n113) );
  AOI22X1 U79 ( .A0(N66), .A1(n125), .B0(N33), .B1(n121), .Y(n112) );
  OAI2BB1X1 U80 ( .A0N(n136), .A1N(\a<20> ), .B0(n133), .Y(n114) );
  NAND2X1 U81 ( .A(n74), .B(n75), .Y(\Result<24> ) );
  AOI22X1 U82 ( .A0(\b<24> ), .A1(n76), .B0(\a<24> ), .B1(n128), .Y(n75) );
  AOI22X1 U83 ( .A0(N70), .A1(n125), .B0(N37), .B1(n124), .Y(n74) );
  OAI2BB1X1 U84 ( .A0N(n136), .A1N(\a<24> ), .B0(n131), .Y(n76) );
  NAND2X1 U85 ( .A(n77), .B(n78), .Y(\Result<23> ) );
  AOI22X1 U86 ( .A0(\b<23> ), .A1(n79), .B0(\a<23> ), .B1(n128), .Y(n78) );
  AOI22X1 U87 ( .A0(N69), .A1(n125), .B0(N36), .B1(n124), .Y(n77) );
  OAI2BB1X1 U88 ( .A0N(n136), .A1N(\a<23> ), .B0(n133), .Y(n79) );
  NAND2X1 U89 ( .A(n28), .B(n29), .Y(\Result<15> ) );
  AOI22X1 U90 ( .A0(\b<15> ), .A1(n30), .B0(\a<15> ), .B1(n128), .Y(n29) );
  AOI22X1 U91 ( .A0(N61), .A1(n126), .B0(N28), .B1(n121), .Y(n28) );
  OAI2BB1X1 U92 ( .A0N(n135), .A1N(\a<15> ), .B0(n129), .Y(n30) );
  NAND2X1 U93 ( .A(n94), .B(n95), .Y(\Result<19> ) );
  AOI22X1 U94 ( .A0(\b<19> ), .A1(n96), .B0(\a<19> ), .B1(n128), .Y(n95) );
  AOI22X1 U95 ( .A0(N65), .A1(n126), .B0(N32), .B1(n121), .Y(n94) );
  OAI2BB1X1 U96 ( .A0N(n136), .A1N(\a<19> ), .B0(n133), .Y(n96) );
  NAND2X1 U97 ( .A(n97), .B(n98), .Y(\Result<18> ) );
  AOI22X1 U98 ( .A0(\b<18> ), .A1(n99), .B0(\a<18> ), .B1(n128), .Y(n98) );
  AOI22X1 U99 ( .A0(N64), .A1(n126), .B0(N31), .B1(n124), .Y(n97) );
  OAI2BB1X1 U100 ( .A0N(n136), .A1N(\a<18> ), .B0(n131), .Y(n99) );
  NAND2X1 U101 ( .A(n100), .B(n101), .Y(\Result<17> ) );
  AOI22X1 U102 ( .A0(\b<17> ), .A1(n102), .B0(\a<17> ), .B1(n19), .Y(n101) );
  AOI22X1 U103 ( .A0(N63), .A1(n126), .B0(N30), .B1(n121), .Y(n100) );
  OAI2BB1X1 U104 ( .A0N(n136), .A1N(\a<17> ), .B0(n133), .Y(n102) );
  NAND2X1 U105 ( .A(n103), .B(n104), .Y(\Result<16> ) );
  AOI22X1 U106 ( .A0(\b<16> ), .A1(n105), .B0(\a<16> ), .B1(n19), .Y(n104) );
  AOI22X1 U107 ( .A0(N62), .A1(n126), .B0(N29), .B1(n121), .Y(n103) );
  OAI2BB1X1 U108 ( .A0N(n136), .A1N(\a<16> ), .B0(n132), .Y(n105) );
  NAND2X1 U109 ( .A(n16), .B(n17), .Y(\Result<11> ) );
  AOI22X1 U110 ( .A0(\b<11> ), .A1(n18), .B0(\a<11> ), .B1(n128), .Y(n17) );
  AOI22X1 U111 ( .A0(N57), .A1(n126), .B0(N24), .B1(n124), .Y(n16) );
  OAI2BB1X1 U112 ( .A0N(n136), .A1N(\a<11> ), .B0(n131), .Y(n18) );
  NAND2X1 U113 ( .A(n22), .B(n23), .Y(\Result<10> ) );
  AOI22X1 U114 ( .A0(\b<10> ), .A1(n24), .B0(\a<10> ), .B1(n128), .Y(n23) );
  AOI22X1 U115 ( .A0(N56), .A1(n126), .B0(N23), .B1(n121), .Y(n22) );
  OAI2BB1X1 U116 ( .A0N(n135), .A1N(\a<10> ), .B0(n131), .Y(n24) );
  NAND2X1 U117 ( .A(n31), .B(n32), .Y(\Result<14> ) );
  AOI22X1 U118 ( .A0(\b<14> ), .A1(n33), .B0(\a<14> ), .B1(n128), .Y(n32) );
  AOI22X1 U119 ( .A0(N60), .A1(n126), .B0(N27), .B1(n121), .Y(n31) );
  OAI2BB1X1 U120 ( .A0N(n135), .A1N(\a<14> ), .B0(n129), .Y(n33) );
  NAND2X1 U121 ( .A(n34), .B(n35), .Y(\Result<13> ) );
  AOI22X1 U122 ( .A0(\b<13> ), .A1(n36), .B0(\a<13> ), .B1(n19), .Y(n35) );
  AOI22X1 U123 ( .A0(N59), .A1(n126), .B0(N26), .B1(n121), .Y(n34) );
  OAI2BB1X1 U124 ( .A0N(n135), .A1N(\a<13> ), .B0(n129), .Y(n36) );
  NAND2X1 U125 ( .A(n37), .B(n38), .Y(\Result<12> ) );
  AOI22X1 U126 ( .A0(\b<12> ), .A1(n39), .B0(\a<12> ), .B1(n128), .Y(n38) );
  AOI22X1 U127 ( .A0(N58), .A1(n126), .B0(N25), .B1(n121), .Y(n37) );
  OAI2BB1X1 U128 ( .A0N(n135), .A1N(\a<12> ), .B0(n130), .Y(n39) );
  NAND2X1 U129 ( .A(n56), .B(n57), .Y(\Result<9> ) );
  AOI22X1 U130 ( .A0(\b<9> ), .A1(n58), .B0(n19), .B1(\a<9> ), .Y(n57) );
  AOI22X1 U131 ( .A0(N55), .A1(n125), .B0(N22), .B1(n121), .Y(n56) );
  OAI2BB1X1 U132 ( .A0N(n136), .A1N(\a<9> ), .B0(n130), .Y(n58) );
  NAND2X1 U133 ( .A(n44), .B(n45), .Y(\Result<5> ) );
  AOI22X1 U134 ( .A0(\b<5> ), .A1(n46), .B0(\a<5> ), .B1(n134), .Y(n45) );
  AOI22X1 U135 ( .A0(N51), .A1(n126), .B0(N18), .B1(n121), .Y(n44) );
  OAI2BB1X1 U136 ( .A0N(n135), .A1N(\a<5> ), .B0(n133), .Y(n46) );
  NAND2X1 U137 ( .A(n47), .B(n48), .Y(\Result<4> ) );
  AOI22X1 U138 ( .A0(\b<4> ), .A1(n49), .B0(\a<4> ), .B1(n128), .Y(n48) );
  AOI22X1 U139 ( .A0(N50), .A1(n125), .B0(N17), .B1(n121), .Y(n47) );
  OAI2BB1X1 U140 ( .A0N(n135), .A1N(\a<4> ), .B0(n132), .Y(n49) );
  NAND2X1 U141 ( .A(n59), .B(n60), .Y(\Result<8> ) );
  AOI22X1 U142 ( .A0(\b<8> ), .A1(n61), .B0(\a<8> ), .B1(n128), .Y(n60) );
  AOI22X1 U143 ( .A0(N54), .A1(n125), .B0(N21), .B1(n124), .Y(n59) );
  OAI2BB1X1 U144 ( .A0N(n136), .A1N(\a<8> ), .B0(n130), .Y(n61) );
  NAND2X1 U145 ( .A(n62), .B(n63), .Y(\Result<7> ) );
  AOI22X1 U146 ( .A0(\b<7> ), .A1(n64), .B0(\a<7> ), .B1(n134), .Y(n63) );
  AOI22X1 U147 ( .A0(N53), .A1(n125), .B0(N20), .B1(n124), .Y(n62) );
  OAI2BB1X1 U148 ( .A0N(n136), .A1N(\a<7> ), .B0(n133), .Y(n64) );
  NAND2X1 U149 ( .A(n65), .B(n66), .Y(\Result<6> ) );
  AOI22X1 U150 ( .A0(\b<6> ), .A1(n67), .B0(\a<6> ), .B1(n128), .Y(n66) );
  AOI22X1 U151 ( .A0(N52), .A1(n125), .B0(N19), .B1(n124), .Y(n65) );
  OAI2BB1X1 U152 ( .A0N(n136), .A1N(\a<6> ), .B0(n131), .Y(n67) );
  NAND2X1 U153 ( .A(n80), .B(n81), .Y(\Result<2> ) );
  AOI22X1 U154 ( .A0(\b<2> ), .A1(n82), .B0(\a<2> ), .B1(n128), .Y(n81) );
  AOI22X1 U155 ( .A0(N48), .A1(n125), .B0(N15), .B1(n124), .Y(n80) );
  OAI2BB1X1 U156 ( .A0N(n136), .A1N(\a<2> ), .B0(n132), .Y(n82) );
  NAND2X1 U157 ( .A(n25), .B(n26), .Y(\Result<0> ) );
  AOI22X1 U158 ( .A0(N46), .A1(n126), .B0(N13), .B1(n121), .Y(n25) );
  NAND2X1 U159 ( .A(n50), .B(n51), .Y(\Result<3> ) );
  AOI22X1 U160 ( .A0(N49), .A1(n125), .B0(N16), .B1(n121), .Y(n50) );
  OAI2BB1X1 U161 ( .A0N(n135), .A1N(n4), .B0(n130), .Y(n52) );
  NAND2X1 U162 ( .A(n115), .B(n116), .Y(\Result<1> ) );
  AOI22X1 U163 ( .A0(N47), .A1(n126), .B0(N14), .B1(n124), .Y(n115) );
  OAI2BB1X1 U164 ( .A0N(n136), .A1N(\a<1> ), .B0(n131), .Y(n117) );
  OAI2BB1X1 U165 ( .A0N(n135), .A1N(n2), .B0(n129), .Y(n27) );
  XOR2X1 U166 ( .A(\b<31> ), .B(\a<31> ), .Y(n120) );
  NOR2BX1 U167 ( .AN(\ALUControl<0> ), .B(n135), .Y(n20) );
  AND2X2 U168 ( .A(\ALUControl<0> ), .B(n135), .Y(n19) );
  OR4X2 U169 ( .A(\Result<12> ), .B(\Result<13> ), .C(\Result<14> ), .D(
        \Result<15> ), .Y(n14) );
  XOR2X1 U170 ( .A(\ALUControl<0> ), .B(n120), .Y(n119) );
  AND2X2 U171 ( .A(N45), .B(n124), .Y(\ALUFlags<1> ) );
  BUFX3 U172 ( .A(\Result<31> ), .Y(\ALUFlags<3> ) );
endmodule


module datapath ( clk, reset, .Adr({\Adr<31> , \Adr<30> , \Adr<29> , \Adr<28> , 
        \Adr<27> , \Adr<26> , \Adr<25> , \Adr<24> , \Adr<23> , \Adr<22> , 
        \Adr<21> , \Adr<20> , \Adr<19> , \Adr<18> , \Adr<17> , \Adr<16> , 
        \Adr<15> , \Adr<14> , \Adr<13> , \Adr<12> , \Adr<11> , \Adr<10> , 
        \Adr<9> , \Adr<8> , \Adr<7> , \Adr<6> , \Adr<5> , \Adr<4> , \Adr<3> , 
        \Adr<2> , \Adr<1> , \Adr<0> }), .WriteData({\WriteData<31> , 
        \WriteData<30> , \WriteData<29> , \WriteData<28> , \WriteData<27> , 
        \WriteData<26> , \WriteData<25> , \WriteData<24> , \WriteData<23> , 
        \WriteData<22> , \WriteData<21> , \WriteData<20> , \WriteData<19> , 
        \WriteData<18> , \WriteData<17> , \WriteData<16> , \WriteData<15> , 
        \WriteData<14> , \WriteData<13> , \WriteData<12> , \WriteData<11> , 
        \WriteData<10> , \WriteData<9> , \WriteData<8> , \WriteData<7> , 
        \WriteData<6> , \WriteData<5> , \WriteData<4> , \WriteData<3> , 
        \WriteData<2> , \WriteData<1> , \WriteData<0> }), .ReadData({
        \ReadData<31> , \ReadData<30> , \ReadData<29> , \ReadData<28> , 
        \ReadData<27> , \ReadData<26> , \ReadData<25> , \ReadData<24> , 
        \ReadData<23> , \ReadData<22> , \ReadData<21> , \ReadData<20> , 
        \ReadData<19> , \ReadData<18> , \ReadData<17> , \ReadData<16> , 
        \ReadData<15> , \ReadData<14> , \ReadData<13> , \ReadData<12> , 
        \ReadData<11> , \ReadData<10> , \ReadData<9> , \ReadData<8> , 
        \ReadData<7> , \ReadData<6> , \ReadData<5> , \ReadData<4> , 
        \ReadData<3> , \ReadData<2> , \ReadData<1> , \ReadData<0> }), .Instr({
        \Instr<31> , \Instr<30> , \Instr<29> , \Instr<28> , \Instr<27> , 
        \Instr<26> , \Instr<25> , \Instr<24> , \Instr<23> , \Instr<22> , 
        \Instr<21> , \Instr<20> , \Instr<19> , \Instr<18> , \Instr<17> , 
        \Instr<16> , \Instr<15> , \Instr<14> , \Instr<13> , \Instr<12> , 
        \Instr<11> , \Instr<10> , \Instr<9> , \Instr<8> , \Instr<7> , 
        \Instr<6> , \Instr<5> , \Instr<4> , \Instr<3> , \Instr<2> , \Instr<1> , 
        \Instr<0> }), .ALUFlags({\ALUFlags<3> , \ALUFlags<2> , \ALUFlags<1> , 
        \ALUFlags<0> }), PCWrite, RegWrite, IRWrite, AdrSrc, .RegSrc({
        \RegSrc<1> , \RegSrc<0> }), .ALUSrcA({\ALUSrcA<1> , \ALUSrcA<0> }), 
    .ALUSrcB({\ALUSrcB<1> , \ALUSrcB<0> }), .ResultSrc({\ResultSrc<1> , 
        \ResultSrc<0> }), .ImmSrc({\ImmSrc<1> , \ImmSrc<0> }), .ALUControl({
        \ALUControl<1> , \ALUControl<0> }) );
  input clk, reset, \ReadData<31> , \ReadData<30> , \ReadData<29> ,
         \ReadData<28> , \ReadData<27> , \ReadData<26> , \ReadData<25> ,
         \ReadData<24> , \ReadData<23> , \ReadData<22> , \ReadData<21> ,
         \ReadData<20> , \ReadData<19> , \ReadData<18> , \ReadData<17> ,
         \ReadData<16> , \ReadData<15> , \ReadData<14> , \ReadData<13> ,
         \ReadData<12> , \ReadData<11> , \ReadData<10> , \ReadData<9> ,
         \ReadData<8> , \ReadData<7> , \ReadData<6> , \ReadData<5> ,
         \ReadData<4> , \ReadData<3> , \ReadData<2> , \ReadData<1> ,
         \ReadData<0> , PCWrite, RegWrite, IRWrite, AdrSrc, \RegSrc<1> ,
         \RegSrc<0> , \ALUSrcA<1> , \ALUSrcA<0> , \ALUSrcB<1> , \ALUSrcB<0> ,
         \ResultSrc<1> , \ResultSrc<0> , \ImmSrc<1> , \ImmSrc<0> ,
         \ALUControl<1> , \ALUControl<0> ;
  output \Adr<31> , \Adr<30> , \Adr<29> , \Adr<28> , \Adr<27> , \Adr<26> ,
         \Adr<25> , \Adr<24> , \Adr<23> , \Adr<22> , \Adr<21> , \Adr<20> ,
         \Adr<19> , \Adr<18> , \Adr<17> , \Adr<16> , \Adr<15> , \Adr<14> ,
         \Adr<13> , \Adr<12> , \Adr<11> , \Adr<10> , \Adr<9> , \Adr<8> ,
         \Adr<7> , \Adr<6> , \Adr<5> , \Adr<4> , \Adr<3> , \Adr<2> , \Adr<1> ,
         \Adr<0> , \WriteData<31> , \WriteData<30> , \WriteData<29> ,
         \WriteData<28> , \WriteData<27> , \WriteData<26> , \WriteData<25> ,
         \WriteData<24> , \WriteData<23> , \WriteData<22> , \WriteData<21> ,
         \WriteData<20> , \WriteData<19> , \WriteData<18> , \WriteData<17> ,
         \WriteData<16> , \WriteData<15> , \WriteData<14> , \WriteData<13> ,
         \WriteData<12> , \WriteData<11> , \WriteData<10> , \WriteData<9> ,
         \WriteData<8> , \WriteData<7> , \WriteData<6> , \WriteData<5> ,
         \WriteData<4> , \WriteData<3> , \WriteData<2> , \WriteData<1> ,
         \WriteData<0> , \Instr<31> , \Instr<30> , \Instr<29> , \Instr<28> ,
         \Instr<27> , \Instr<26> , \Instr<25> , \Instr<24> , \Instr<23> ,
         \Instr<22> , \Instr<21> , \Instr<20> , \Instr<19> , \Instr<18> ,
         \Instr<17> , \Instr<16> , \Instr<15> , \Instr<14> , \Instr<13> ,
         \Instr<12> , \Instr<11> , \Instr<10> , \Instr<9> , \Instr<8> ,
         \Instr<7> , \Instr<6> , \Instr<5> , \Instr<4> , \Instr<3> ,
         \Instr<2> , \Instr<1> , \Instr<0> , \ALUFlags<3> , \ALUFlags<2> ,
         \ALUFlags<1> , \ALUFlags<0> ;
  wire   \PC<31> , \PC<30> , \PC<29> , \PC<28> , \PC<27> , \PC<26> , \PC<25> ,
         \PC<24> , \PC<23> , \PC<22> , \PC<21> , \PC<20> , \PC<19> , \PC<18> ,
         \PC<17> , \PC<16> , \PC<15> , \PC<14> , \PC<13> , \PC<12> , \PC<11> ,
         \PC<10> , \PC<9> , \PC<8> , \PC<7> , \PC<6> , \PC<5> , \PC<4> ,
         \PC<3> , \PC<2> , \PC<1> , \PC<0> , \Data<31> , \Data<30> ,
         \Data<29> , \Data<28> , \Data<27> , \Data<26> , \Data<25> ,
         \Data<24> , \Data<23> , \Data<22> , \Data<21> , \Data<20> ,
         \Data<19> , \Data<18> , \Data<17> , \Data<16> , \Data<15> ,
         \Data<14> , \Data<13> , \Data<12> , \Data<11> , \Data<10> , \Data<9> ,
         \Data<8> , \Data<7> , \Data<6> , \Data<5> , \Data<4> , \Data<3> ,
         \Data<2> , \Data<1> , \Data<0> , \RD1<31> , \RD1<30> , \RD1<29> ,
         \RD1<28> , \RD1<27> , \RD1<26> , \RD1<25> , \RD1<24> , \RD1<23> ,
         \RD1<22> , \RD1<21> , \RD1<20> , \RD1<19> , \RD1<18> , \RD1<17> ,
         \RD1<16> , \RD1<15> , \RD1<14> , \RD1<13> , \RD1<12> , \RD1<11> ,
         \RD1<10> , \RD1<9> , \RD1<8> , \RD1<7> , \RD1<6> , \RD1<5> , \RD1<4> ,
         \RD1<3> , \RD1<2> , \RD1<1> , \RD1<0> , \A<31> , \A<30> , \A<29> ,
         \A<28> , \A<27> , \A<26> , \A<25> , \A<24> , \A<23> , \A<22> ,
         \A<21> , \A<20> , \A<19> , \A<18> , \A<17> , \A<16> , \A<15> ,
         \A<14> , \A<13> , \A<12> , \A<11> , \A<10> , \A<9> , \A<8> , \A<7> ,
         \A<6> , \A<5> , \A<4> , \A<3> , \A<2> , \A<1> , \A<0> , \RD2<31> ,
         \RD2<30> , \RD2<29> , \RD2<28> , \RD2<27> , \RD2<26> , \RD2<25> ,
         \RD2<24> , \RD2<23> , \RD2<22> , \RD2<21> , \RD2<20> , \RD2<19> ,
         \RD2<18> , \RD2<17> , \RD2<16> , \RD2<15> , \RD2<14> , \RD2<13> ,
         \RD2<12> , \RD2<11> , \RD2<10> , \RD2<9> , \RD2<8> , \RD2<7> ,
         \RD2<6> , \RD2<5> , \RD2<4> , \RD2<3> , \RD2<2> , \RD2<1> , \RD2<0> ,
         \ALUResult<31> , \ALUResult<30> , \ALUResult<29> , \ALUResult<28> ,
         \ALUResult<27> , \ALUResult<26> , \ALUResult<25> , \ALUResult<24> ,
         \ALUResult<23> , \ALUResult<22> , \ALUResult<21> , \ALUResult<20> ,
         \ALUResult<19> , \ALUResult<18> , \ALUResult<17> , \ALUResult<16> ,
         \ALUResult<15> , \ALUResult<14> , \ALUResult<13> , \ALUResult<12> ,
         \ALUResult<11> , \ALUResult<10> , \ALUResult<9> , \ALUResult<8> ,
         \ALUResult<7> , \ALUResult<6> , \ALUResult<5> , \ALUResult<4> ,
         \ALUResult<3> , \ALUResult<2> , \ALUResult<1> , \ALUResult<0> ,
         \ALUOut<31> , \ALUOut<30> , \ALUOut<29> , \ALUOut<28> , \ALUOut<27> ,
         \ALUOut<26> , \ALUOut<25> , \ALUOut<24> , \ALUOut<23> , \ALUOut<22> ,
         \ALUOut<21> , \ALUOut<20> , \ALUOut<19> , \ALUOut<18> , \ALUOut<17> ,
         \ALUOut<16> , \ALUOut<15> , \ALUOut<14> , \ALUOut<13> , \ALUOut<12> ,
         \ALUOut<11> , \ALUOut<10> , \ALUOut<9> , \ALUOut<8> , \ALUOut<7> ,
         \ALUOut<6> , \ALUOut<5> , \ALUOut<4> , \ALUOut<3> , \ALUOut<2> ,
         \ALUOut<1> , \ALUOut<0> , \Result<31> , \Result<30> , \Result<29> ,
         \Result<28> , \Result<27> , \Result<26> , \Result<25> , \Result<24> ,
         \Result<23> , \Result<22> , \Result<21> , \Result<20> , \Result<19> ,
         \Result<18> , \Result<17> , \Result<16> , \Result<15> , \Result<14> ,
         \Result<13> , \Result<12> , \Result<11> , \Result<10> , \Result<9> ,
         \Result<8> , \Result<7> , \Result<6> , \Result<5> , \Result<4> ,
         \Result<3> , \Result<2> , \Result<1> , \Result<0> , \RA1<3> ,
         \RA1<2> , \RA1<1> , \RA1<0> , \RA2<3> , \RA2<2> , \RA2<1> , \RA2<0> ,
         \SrcA<31> , \SrcA<30> , \SrcA<29> , \SrcA<28> , \SrcA<27> ,
         \SrcA<26> , \SrcA<25> , \SrcA<24> , \SrcA<23> , \SrcA<22> ,
         \SrcA<21> , \SrcA<20> , \SrcA<19> , \SrcA<18> , \SrcA<17> ,
         \SrcA<16> , \SrcA<15> , \SrcA<14> , \SrcA<13> , \SrcA<12> ,
         \SrcA<11> , \SrcA<10> , \SrcA<9> , \SrcA<8> , \SrcA<7> , \SrcA<6> ,
         \SrcA<5> , \SrcA<4> , \SrcA<3> , \SrcA<2> , \SrcA<1> , \SrcA<0> ,
         \ExtImm<31> , \ExtImm<30> , \ExtImm<29> , \ExtImm<28> , \ExtImm<27> ,
         \ExtImm<26> , \ExtImm<25> , \ExtImm<24> , \ExtImm<23> , \ExtImm<22> ,
         \ExtImm<21> , \ExtImm<20> , \ExtImm<19> , \ExtImm<18> , \ExtImm<17> ,
         \ExtImm<16> , \ExtImm<15> , \ExtImm<14> , \ExtImm<13> , \ExtImm<12> ,
         \ExtImm<11> , \ExtImm<10> , \ExtImm<9> , \ExtImm<8> , \ExtImm<7> ,
         \ExtImm<6> , \ExtImm<5> , \ExtImm<4> , \ExtImm<3> , \ExtImm<2> ,
         \ExtImm<1> , \ExtImm<0> , \SrcB<31> , \SrcB<30> , \SrcB<29> ,
         \SrcB<28> , \SrcB<27> , \SrcB<26> , \SrcB<25> , \SrcB<24> ,
         \SrcB<23> , \SrcB<22> , \SrcB<21> , \SrcB<20> , \SrcB<19> ,
         \SrcB<18> , \SrcB<17> , \SrcB<16> , \SrcB<15> , \SrcB<14> ,
         \SrcB<13> , \SrcB<12> , \SrcB<11> , \SrcB<10> , \SrcB<9> , \SrcB<8> ,
         \SrcB<7> , \SrcB<6> , \SrcB<5> , \SrcB<4> , \SrcB<3> , \SrcB<2> ,
         \SrcB<1> , \SrcB<0> , n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11,
         n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25,
         n26, n27, n28, n29, n30, n31, n32, n33, n34;

  flopenr_WIDTH32_0 pcreg ( .clk(clk), .reset(reset), .en(n33), .d({n2, n1, 
        \Result<29> , \Result<28> , \Result<27> , \Result<26> , \Result<25> , 
        \Result<24> , \Result<23> , \Result<22> , \Result<21> , \Result<20> , 
        \Result<19> , \Result<18> , \Result<17> , \Result<16> , \Result<15> , 
        \Result<14> , \Result<13> , \Result<12> , \Result<11> , \Result<10> , 
        \Result<9> , \Result<8> , \Result<7> , \Result<6> , \Result<5> , 
        \Result<4> , \Result<3> , \Result<2> , \Result<1> , \Result<0> }), .q(
        {\PC<31> , \PC<30> , \PC<29> , \PC<28> , \PC<27> , \PC<26> , \PC<25> , 
        \PC<24> , \PC<23> , \PC<22> , \PC<21> , \PC<20> , \PC<19> , \PC<18> , 
        \PC<17> , \PC<16> , \PC<15> , \PC<14> , \PC<13> , \PC<12> , \PC<11> , 
        \PC<10> , \PC<9> , \PC<8> , \PC<7> , \PC<6> , \PC<5> , \PC<4> , 
        \PC<3> , \PC<2> , \PC<1> , \PC<0> }) );
  flopenr_WIDTH32_1 instrreg ( .clk(clk), .reset(reset), .en(n31), .d({
        \ReadData<31> , \ReadData<30> , \ReadData<29> , \ReadData<28> , 
        \ReadData<27> , \ReadData<26> , \ReadData<25> , \ReadData<24> , 
        \ReadData<23> , \ReadData<22> , \ReadData<21> , \ReadData<20> , 
        \ReadData<19> , \ReadData<18> , \ReadData<17> , \ReadData<16> , 
        \ReadData<15> , \ReadData<14> , \ReadData<13> , \ReadData<12> , 
        \ReadData<11> , \ReadData<10> , \ReadData<9> , \ReadData<8> , 
        \ReadData<7> , \ReadData<6> , \ReadData<5> , \ReadData<4> , 
        \ReadData<3> , \ReadData<2> , \ReadData<1> , \ReadData<0> }), .q({
        \Instr<31> , \Instr<30> , \Instr<29> , \Instr<28> , \Instr<27> , 
        \Instr<26> , \Instr<25> , \Instr<24> , \Instr<23> , \Instr<22> , 
        \Instr<21> , \Instr<20> , \Instr<19> , \Instr<18> , \Instr<17> , 
        \Instr<16> , \Instr<15> , \Instr<14> , \Instr<13> , \Instr<12> , 
        \Instr<11> , \Instr<10> , \Instr<9> , \Instr<8> , \Instr<7> , 
        \Instr<6> , \Instr<5> , \Instr<4> , \Instr<3> , \Instr<2> , \Instr<1> , 
        \Instr<0> }) );
  flopr_WIDTH32_0 datareg ( .clk(clk), .reset(reset), .d({\ReadData<31> , 
        \ReadData<30> , \ReadData<29> , \ReadData<28> , \ReadData<27> , 
        \ReadData<26> , \ReadData<25> , \ReadData<24> , \ReadData<23> , 
        \ReadData<22> , \ReadData<21> , \ReadData<20> , \ReadData<19> , 
        \ReadData<18> , \ReadData<17> , \ReadData<16> , \ReadData<15> , 
        \ReadData<14> , \ReadData<13> , \ReadData<12> , \ReadData<11> , 
        \ReadData<10> , \ReadData<9> , \ReadData<8> , \ReadData<7> , 
        \ReadData<6> , \ReadData<5> , \ReadData<4> , \ReadData<3> , 
        \ReadData<2> , \ReadData<1> , \ReadData<0> }), .q({\Data<31> , 
        \Data<30> , \Data<29> , \Data<28> , \Data<27> , \Data<26> , \Data<25> , 
        \Data<24> , \Data<23> , \Data<22> , \Data<21> , \Data<20> , \Data<19> , 
        \Data<18> , \Data<17> , \Data<16> , \Data<15> , \Data<14> , \Data<13> , 
        \Data<12> , \Data<11> , \Data<10> , \Data<9> , \Data<8> , \Data<7> , 
        \Data<6> , \Data<5> , \Data<4> , \Data<3> , \Data<2> , \Data<1> , 
        \Data<0> }) );
  flopr_WIDTH32_3 rd1reg ( .clk(clk), .reset(reset), .d({\RD1<31> , \RD1<30> , 
        \RD1<29> , \RD1<28> , \RD1<27> , \RD1<26> , \RD1<25> , \RD1<24> , 
        \RD1<23> , \RD1<22> , \RD1<21> , \RD1<20> , \RD1<19> , \RD1<18> , 
        \RD1<17> , \RD1<16> , \RD1<15> , \RD1<14> , \RD1<13> , \RD1<12> , 
        \RD1<11> , \RD1<10> , \RD1<9> , \RD1<8> , \RD1<7> , \RD1<6> , \RD1<5> , 
        \RD1<4> , \RD1<3> , \RD1<2> , \RD1<1> , \RD1<0> }), .q({\A<31> , 
        \A<30> , \A<29> , \A<28> , \A<27> , \A<26> , \A<25> , \A<24> , \A<23> , 
        \A<22> , \A<21> , \A<20> , \A<19> , \A<18> , \A<17> , \A<16> , \A<15> , 
        \A<14> , \A<13> , \A<12> , \A<11> , \A<10> , \A<9> , \A<8> , \A<7> , 
        \A<6> , \A<5> , \A<4> , \A<3> , \A<2> , \A<1> , \A<0> }) );
  flopr_WIDTH32_2 rd2reg ( .clk(clk), .reset(reset), .d({\RD2<31> , \RD2<30> , 
        \RD2<29> , \RD2<28> , \RD2<27> , \RD2<26> , \RD2<25> , \RD2<24> , 
        \RD2<23> , \RD2<22> , \RD2<21> , \RD2<20> , \RD2<19> , \RD2<18> , 
        \RD2<17> , \RD2<16> , \RD2<15> , \RD2<14> , \RD2<13> , \RD2<12> , 
        \RD2<11> , \RD2<10> , \RD2<9> , \RD2<8> , \RD2<7> , \RD2<6> , \RD2<5> , 
        \RD2<4> , \RD2<3> , \RD2<2> , \RD2<1> , \RD2<0> }), .q({
        \WriteData<31> , \WriteData<30> , \WriteData<29> , \WriteData<28> , 
        \WriteData<27> , \WriteData<26> , \WriteData<25> , \WriteData<24> , 
        \WriteData<23> , \WriteData<22> , \WriteData<21> , \WriteData<20> , 
        \WriteData<19> , \WriteData<18> , \WriteData<17> , \WriteData<16> , 
        \WriteData<15> , \WriteData<14> , \WriteData<13> , \WriteData<12> , 
        \WriteData<11> , \WriteData<10> , \WriteData<9> , \WriteData<8> , 
        \WriteData<7> , \WriteData<6> , \WriteData<5> , \WriteData<4> , 
        \WriteData<3> , \WriteData<2> , \WriteData<1> , \WriteData<0> }) );
  flopr_WIDTH32_1 alureg ( .clk(clk), .reset(reset), .d({\ALUResult<31> , 
        \ALUResult<30> , \ALUResult<29> , \ALUResult<28> , \ALUResult<27> , 
        \ALUResult<26> , \ALUResult<25> , \ALUResult<24> , \ALUResult<23> , 
        \ALUResult<22> , \ALUResult<21> , \ALUResult<20> , \ALUResult<19> , 
        \ALUResult<18> , \ALUResult<17> , \ALUResult<16> , \ALUResult<15> , 
        \ALUResult<14> , \ALUResult<13> , \ALUResult<12> , \ALUResult<11> , 
        \ALUResult<10> , \ALUResult<9> , \ALUResult<8> , \ALUResult<7> , 
        \ALUResult<6> , \ALUResult<5> , \ALUResult<4> , \ALUResult<3> , 
        \ALUResult<2> , \ALUResult<1> , \ALUResult<0> }), .q({\ALUOut<31> , 
        \ALUOut<30> , \ALUOut<29> , \ALUOut<28> , \ALUOut<27> , \ALUOut<26> , 
        \ALUOut<25> , \ALUOut<24> , \ALUOut<23> , \ALUOut<22> , \ALUOut<21> , 
        \ALUOut<20> , \ALUOut<19> , \ALUOut<18> , \ALUOut<17> , \ALUOut<16> , 
        \ALUOut<15> , \ALUOut<14> , \ALUOut<13> , \ALUOut<12> , \ALUOut<11> , 
        \ALUOut<10> , \ALUOut<9> , \ALUOut<8> , \ALUOut<7> , \ALUOut<6> , 
        \ALUOut<5> , \ALUOut<4> , \ALUOut<3> , \ALUOut<2> , \ALUOut<1> , 
        \ALUOut<0> }) );
  mux2_WIDTH32 adrmux ( .d0({\PC<31> , \PC<30> , \PC<29> , \PC<28> , \PC<27> , 
        \PC<26> , \PC<25> , \PC<24> , \PC<23> , \PC<22> , \PC<21> , \PC<20> , 
        \PC<19> , \PC<18> , \PC<17> , \PC<16> , \PC<15> , \PC<14> , \PC<13> , 
        \PC<12> , \PC<11> , \PC<10> , \PC<9> , \PC<8> , \PC<7> , \PC<6> , 
        \PC<5> , \PC<4> , \PC<3> , \PC<2> , \PC<1> , \PC<0> }), .d1({n2, n1, 
        \Result<29> , \Result<28> , \Result<27> , \Result<26> , \Result<25> , 
        \Result<24> , \Result<23> , \Result<22> , \Result<21> , \Result<20> , 
        \Result<19> , \Result<18> , \Result<17> , \Result<16> , \Result<15> , 
        \Result<14> , \Result<13> , \Result<12> , \Result<11> , \Result<10> , 
        \Result<9> , \Result<8> , \Result<7> , \Result<6> , \Result<5> , 
        \Result<4> , \Result<3> , \Result<2> , \Result<1> , \Result<0> }), .s(
        n29), .y({\Adr<31> , \Adr<30> , \Adr<29> , \Adr<28> , \Adr<27> , 
        \Adr<26> , \Adr<25> , \Adr<24> , \Adr<23> , \Adr<22> , \Adr<21> , 
        \Adr<20> , \Adr<19> , \Adr<18> , \Adr<17> , \Adr<16> , \Adr<15> , 
        \Adr<14> , \Adr<13> , \Adr<12> , \Adr<11> , \Adr<10> , \Adr<9> , 
        \Adr<8> , \Adr<7> , \Adr<6> , \Adr<5> , \Adr<4> , \Adr<3> , \Adr<2> , 
        \Adr<1> , \Adr<0> }) );
  mux2_WIDTH4_0 ra1mux ( .d0({\Instr<19> , \Instr<18> , \Instr<17> , 
        \Instr<16> }), .d1({1'b1, 1'b1, 1'b1, 1'b1}), .s(\RegSrc<0> ), .y({
        \RA1<3> , \RA1<2> , \RA1<1> , \RA1<0> }) );
  mux2_WIDTH4_1 ra2mux ( .d0({\Instr<3> , \Instr<2> , \Instr<1> , \Instr<0> }), 
        .d1({\Instr<15> , \Instr<14> , \Instr<13> , \Instr<12> }), .s(
        \RegSrc<1> ), .y({\RA2<3> , \RA2<2> , \RA2<1> , \RA2<0> }) );
  mux3_WIDTH32_0 srcAmux ( .d0({\A<31> , \A<30> , \A<29> , \A<28> , \A<27> , 
        \A<26> , \A<25> , \A<24> , \A<23> , \A<22> , \A<21> , \A<20> , \A<19> , 
        \A<18> , \A<17> , \A<16> , \A<15> , \A<14> , \A<13> , \A<12> , \A<11> , 
        \A<10> , \A<9> , \A<8> , \A<7> , \A<6> , \A<5> , \A<4> , \A<3> , 
        \A<2> , \A<1> , \A<0> }), .d1({\PC<31> , \PC<30> , \PC<29> , \PC<28> , 
        \PC<27> , \PC<26> , \PC<25> , \PC<24> , \PC<23> , \PC<22> , \PC<21> , 
        \PC<20> , \PC<19> , \PC<18> , \PC<17> , \PC<16> , \PC<15> , \PC<14> , 
        \PC<13> , \PC<12> , \PC<11> , \PC<10> , \PC<9> , \PC<8> , \PC<7> , 
        \PC<6> , \PC<5> , \PC<4> , \PC<3> , \PC<2> , \PC<1> , \PC<0> }), .d2({
        \ALUOut<31> , \ALUOut<30> , \ALUOut<29> , \ALUOut<28> , \ALUOut<27> , 
        \ALUOut<26> , \ALUOut<25> , \ALUOut<24> , \ALUOut<23> , \ALUOut<22> , 
        \ALUOut<21> , \ALUOut<20> , \ALUOut<19> , \ALUOut<18> , \ALUOut<17> , 
        \ALUOut<16> , \ALUOut<15> , \ALUOut<14> , \ALUOut<13> , \ALUOut<12> , 
        \ALUOut<11> , \ALUOut<10> , \ALUOut<9> , \ALUOut<8> , \ALUOut<7> , 
        \ALUOut<6> , \ALUOut<5> , \ALUOut<4> , \ALUOut<3> , \ALUOut<2> , 
        \ALUOut<1> , \ALUOut<0> }), .s({n27, n25}), .y({\SrcA<31> , \SrcA<30> , 
        \SrcA<29> , \SrcA<28> , \SrcA<27> , \SrcA<26> , \SrcA<25> , \SrcA<24> , 
        \SrcA<23> , \SrcA<22> , \SrcA<21> , \SrcA<20> , \SrcA<19> , \SrcA<18> , 
        \SrcA<17> , \SrcA<16> , \SrcA<15> , \SrcA<14> , \SrcA<13> , \SrcA<12> , 
        \SrcA<11> , \SrcA<10> , \SrcA<9> , \SrcA<8> , \SrcA<7> , \SrcA<6> , 
        \SrcA<5> , \SrcA<4> , \SrcA<3> , \SrcA<2> , \SrcA<1> , \SrcA<0> }) );
  mux3_WIDTH32_2 srcBmux ( .d0({\WriteData<31> , \WriteData<30> , 
        \WriteData<29> , \WriteData<28> , \WriteData<27> , \WriteData<26> , 
        \WriteData<25> , \WriteData<24> , \WriteData<23> , \WriteData<22> , 
        \WriteData<21> , \WriteData<20> , \WriteData<19> , \WriteData<18> , 
        \WriteData<17> , \WriteData<16> , \WriteData<15> , \WriteData<14> , 
        \WriteData<13> , \WriteData<12> , \WriteData<11> , \WriteData<10> , 
        \WriteData<9> , \WriteData<8> , \WriteData<7> , \WriteData<6> , 
        \WriteData<5> , \WriteData<4> , \WriteData<3> , \WriteData<2> , 
        \WriteData<1> , \WriteData<0> }), .d1({\ExtImm<31> , \ExtImm<30> , 
        \ExtImm<29> , \ExtImm<28> , \ExtImm<27> , \ExtImm<26> , \ExtImm<25> , 
        \ExtImm<24> , \ExtImm<23> , \ExtImm<22> , \ExtImm<21> , \ExtImm<20> , 
        \ExtImm<19> , \ExtImm<18> , \ExtImm<17> , \ExtImm<16> , \ExtImm<15> , 
        \ExtImm<14> , \ExtImm<13> , \ExtImm<12> , \ExtImm<11> , \ExtImm<10> , 
        \ExtImm<9> , \ExtImm<8> , \ExtImm<7> , \ExtImm<6> , \ExtImm<5> , 
        \ExtImm<4> , \ExtImm<3> , \ExtImm<2> , \ExtImm<1> , \ExtImm<0> }), 
        .d2({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0}), .s({n23, 
        \ALUSrcB<0> }), .y({\SrcB<31> , \SrcB<30> , \SrcB<29> , \SrcB<28> , 
        \SrcB<27> , \SrcB<26> , \SrcB<25> , \SrcB<24> , \SrcB<23> , \SrcB<22> , 
        \SrcB<21> , \SrcB<20> , \SrcB<19> , \SrcB<18> , \SrcB<17> , \SrcB<16> , 
        \SrcB<15> , \SrcB<14> , \SrcB<13> , \SrcB<12> , \SrcB<11> , \SrcB<10> , 
        \SrcB<9> , \SrcB<8> , \SrcB<7> , \SrcB<6> , \SrcB<5> , \SrcB<4> , 
        \SrcB<3> , \SrcB<2> , \SrcB<1> , \SrcB<0> }) );
  mux3_WIDTH32_1 alumux ( .d0({\ALUOut<31> , \ALUOut<30> , \ALUOut<29> , 
        \ALUOut<28> , \ALUOut<27> , \ALUOut<26> , \ALUOut<25> , \ALUOut<24> , 
        \ALUOut<23> , \ALUOut<22> , \ALUOut<21> , \ALUOut<20> , \ALUOut<19> , 
        \ALUOut<18> , \ALUOut<17> , \ALUOut<16> , \ALUOut<15> , \ALUOut<14> , 
        \ALUOut<13> , \ALUOut<12> , \ALUOut<11> , \ALUOut<10> , \ALUOut<9> , 
        \ALUOut<8> , \ALUOut<7> , \ALUOut<6> , \ALUOut<5> , \ALUOut<4> , 
        \ALUOut<3> , \ALUOut<2> , \ALUOut<1> , \ALUOut<0> }), .d1({\Data<31> , 
        \Data<30> , \Data<29> , \Data<28> , \Data<27> , \Data<26> , \Data<25> , 
        \Data<24> , \Data<23> , \Data<22> , \Data<21> , \Data<20> , \Data<19> , 
        \Data<18> , \Data<17> , \Data<16> , \Data<15> , \Data<14> , \Data<13> , 
        \Data<12> , \Data<11> , \Data<10> , \Data<9> , \Data<8> , \Data<7> , 
        \Data<6> , \Data<5> , \Data<4> , \Data<3> , \Data<2> , \Data<1> , 
        \Data<0> }), .d2({\ALUResult<31> , \ALUResult<30> , \ALUResult<29> , 
        \ALUResult<28> , \ALUResult<27> , \ALUResult<26> , \ALUResult<25> , 
        \ALUResult<24> , \ALUResult<23> , \ALUResult<22> , \ALUResult<21> , 
        \ALUResult<20> , \ALUResult<19> , \ALUResult<18> , \ALUResult<17> , 
        \ALUResult<16> , \ALUResult<15> , \ALUResult<14> , \ALUResult<13> , 
        \ALUResult<12> , \ALUResult<11> , \ALUResult<10> , \ALUResult<9> , 
        \ALUResult<8> , \ALUResult<7> , \ALUResult<6> , \ALUResult<5> , 
        \ALUResult<4> , \ALUResult<3> , \ALUResult<2> , \ALUResult<1> , 
        \ALUResult<0> }), .s({n21, \ResultSrc<0> }), .y({\Result<31> , 
        \Result<30> , \Result<29> , \Result<28> , \Result<27> , \Result<26> , 
        \Result<25> , \Result<24> , \Result<23> , \Result<22> , \Result<21> , 
        \Result<20> , \Result<19> , \Result<18> , \Result<17> , \Result<16> , 
        \Result<15> , \Result<14> , \Result<13> , \Result<12> , \Result<11> , 
        \Result<10> , \Result<9> , \Result<8> , \Result<7> , \Result<6> , 
        \Result<5> , \Result<4> , \Result<3> , \Result<2> , \Result<1> , 
        \Result<0> }) );
  regfile rf ( .clk(clk), .we3(RegWrite), .ra1({n17, n15, n13, n11}), .ra2({n9, 
        n7, n5, n3}), .wa3({\Instr<15> , \Instr<14> , \Instr<13> , \Instr<12> }), .wd3({n2, n1, \Result<29> , \Result<28> , \Result<27> , \Result<26> , 
        \Result<25> , \Result<24> , \Result<23> , \Result<22> , \Result<21> , 
        \Result<20> , \Result<19> , \Result<18> , \Result<17> , \Result<16> , 
        \Result<15> , \Result<14> , \Result<13> , \Result<12> , \Result<11> , 
        \Result<10> , \Result<9> , \Result<8> , \Result<7> , \Result<6> , 
        \Result<5> , \Result<4> , \Result<3> , \Result<2> , \Result<1> , 
        \Result<0> }), .r15({n2, n1, \Result<29> , \Result<28> , \Result<27> , 
        \Result<26> , \Result<25> , \Result<24> , \Result<23> , \Result<22> , 
        \Result<21> , \Result<20> , \Result<19> , \Result<18> , \Result<17> , 
        \Result<16> , \Result<15> , \Result<14> , \Result<13> , \Result<12> , 
        \Result<11> , \Result<10> , \Result<9> , \Result<8> , \Result<7> , 
        \Result<6> , \Result<5> , \Result<4> , \Result<3> , \Result<2> , 
        \Result<1> , \Result<0> }), .rd1({\RD1<31> , \RD1<30> , \RD1<29> , 
        \RD1<28> , \RD1<27> , \RD1<26> , \RD1<25> , \RD1<24> , \RD1<23> , 
        \RD1<22> , \RD1<21> , \RD1<20> , \RD1<19> , \RD1<18> , \RD1<17> , 
        \RD1<16> , \RD1<15> , \RD1<14> , \RD1<13> , \RD1<12> , \RD1<11> , 
        \RD1<10> , \RD1<9> , \RD1<8> , \RD1<7> , \RD1<6> , \RD1<5> , \RD1<4> , 
        \RD1<3> , \RD1<2> , \RD1<1> , \RD1<0> }), .rd2({\RD2<31> , \RD2<30> , 
        \RD2<29> , \RD2<28> , \RD2<27> , \RD2<26> , \RD2<25> , \RD2<24> , 
        \RD2<23> , \RD2<22> , \RD2<21> , \RD2<20> , \RD2<19> , \RD2<18> , 
        \RD2<17> , \RD2<16> , \RD2<15> , \RD2<14> , \RD2<13> , \RD2<12> , 
        \RD2<11> , \RD2<10> , \RD2<9> , \RD2<8> , \RD2<7> , \RD2<6> , \RD2<5> , 
        \RD2<4> , \RD2<3> , \RD2<2> , \RD2<1> , \RD2<0> }) );
  extend ext ( .Instr({\Instr<23> , \Instr<22> , \Instr<21> , \Instr<20> , 
        \Instr<19> , \Instr<18> , \Instr<17> , \Instr<16> , \Instr<15> , 
        \Instr<14> , \Instr<13> , \Instr<12> , \Instr<11> , \Instr<10> , 
        \Instr<9> , \Instr<8> , \Instr<7> , \Instr<6> , \Instr<5> , \Instr<4> , 
        \Instr<3> , \Instr<2> , \Instr<1> , \Instr<0> }), .ImmSrc({\ImmSrc<1> , 
        \ImmSrc<0> }), .ExtImm({\ExtImm<31> , \ExtImm<30> , \ExtImm<29> , 
        \ExtImm<28> , \ExtImm<27> , \ExtImm<26> , \ExtImm<25> , \ExtImm<24> , 
        \ExtImm<23> , \ExtImm<22> , \ExtImm<21> , \ExtImm<20> , \ExtImm<19> , 
        \ExtImm<18> , \ExtImm<17> , \ExtImm<16> , \ExtImm<15> , \ExtImm<14> , 
        \ExtImm<13> , \ExtImm<12> , \ExtImm<11> , \ExtImm<10> , \ExtImm<9> , 
        \ExtImm<8> , \ExtImm<7> , \ExtImm<6> , \ExtImm<5> , \ExtImm<4> , 
        \ExtImm<3> , \ExtImm<2> , \ExtImm<1> , \ExtImm<0> }) );
  alu alu ( .a({\SrcA<31> , \SrcA<30> , \SrcA<29> , \SrcA<28> , \SrcA<27> , 
        \SrcA<26> , \SrcA<25> , \SrcA<24> , \SrcA<23> , \SrcA<22> , \SrcA<21> , 
        \SrcA<20> , \SrcA<19> , \SrcA<18> , \SrcA<17> , \SrcA<16> , \SrcA<15> , 
        \SrcA<14> , \SrcA<13> , \SrcA<12> , \SrcA<11> , \SrcA<10> , \SrcA<9> , 
        \SrcA<8> , \SrcA<7> , \SrcA<6> , \SrcA<5> , \SrcA<4> , \SrcA<3> , 
        \SrcA<2> , \SrcA<1> , \SrcA<0> }), .b({\SrcB<31> , \SrcB<30> , 
        \SrcB<29> , \SrcB<28> , \SrcB<27> , \SrcB<26> , \SrcB<25> , \SrcB<24> , 
        \SrcB<23> , \SrcB<22> , \SrcB<21> , \SrcB<20> , \SrcB<19> , \SrcB<18> , 
        \SrcB<17> , \SrcB<16> , \SrcB<15> , \SrcB<14> , \SrcB<13> , \SrcB<12> , 
        \SrcB<11> , \SrcB<10> , \SrcB<9> , \SrcB<8> , \SrcB<7> , \SrcB<6> , 
        \SrcB<5> , \SrcB<4> , \SrcB<3> , \SrcB<2> , \SrcB<1> , \SrcB<0> }), 
        .ALUControl({n19, \ALUControl<0> }), .Result({\ALUResult<31> , 
        \ALUResult<30> , \ALUResult<29> , \ALUResult<28> , \ALUResult<27> , 
        \ALUResult<26> , \ALUResult<25> , \ALUResult<24> , \ALUResult<23> , 
        \ALUResult<22> , \ALUResult<21> , \ALUResult<20> , \ALUResult<19> , 
        \ALUResult<18> , \ALUResult<17> , \ALUResult<16> , \ALUResult<15> , 
        \ALUResult<14> , \ALUResult<13> , \ALUResult<12> , \ALUResult<11> , 
        \ALUResult<10> , \ALUResult<9> , \ALUResult<8> , \ALUResult<7> , 
        \ALUResult<6> , \ALUResult<5> , \ALUResult<4> , \ALUResult<3> , 
        \ALUResult<2> , \ALUResult<1> , \ALUResult<0> }), .ALUFlags({
        \ALUFlags<3> , \ALUFlags<2> , \ALUFlags<1> , \ALUFlags<0> }) );
  BUFX12 U3 ( .A(\Result<30> ), .Y(n1) );
  BUFX20 U4 ( .A(\Result<31> ), .Y(n2) );
  INVX4 U5 ( .A(n24), .Y(n23) );
  INVX1 U6 ( .A(n26), .Y(n25) );
  INVX1 U7 ( .A(\ALUSrcA<0> ), .Y(n26) );
  INVX1 U8 ( .A(n28), .Y(n27) );
  INVX4 U9 ( .A(\ALUSrcA<1> ), .Y(n28) );
  INVX1 U10 ( .A(\ALUSrcB<1> ), .Y(n24) );
  INVX1 U11 ( .A(n22), .Y(n21) );
  INVX1 U12 ( .A(\ResultSrc<1> ), .Y(n22) );
  INVX1 U13 ( .A(n32), .Y(n31) );
  INVX1 U14 ( .A(IRWrite), .Y(n32) );
  INVX1 U15 ( .A(n34), .Y(n33) );
  INVX1 U16 ( .A(PCWrite), .Y(n34) );
  INVX1 U17 ( .A(n20), .Y(n19) );
  INVX1 U18 ( .A(\ALUControl<1> ), .Y(n20) );
  INVX1 U19 ( .A(n30), .Y(n29) );
  INVX1 U20 ( .A(AdrSrc), .Y(n30) );
  INVX1 U21 ( .A(n12), .Y(n11) );
  INVX1 U22 ( .A(\RA1<0> ), .Y(n12) );
  INVX1 U23 ( .A(n4), .Y(n3) );
  INVX1 U24 ( .A(\RA2<0> ), .Y(n4) );
  INVX1 U25 ( .A(n10), .Y(n9) );
  INVX1 U26 ( .A(\RA2<3> ), .Y(n10) );
  INVX1 U27 ( .A(n14), .Y(n13) );
  INVX1 U28 ( .A(\RA1<1> ), .Y(n14) );
  INVX1 U29 ( .A(n6), .Y(n5) );
  INVX1 U30 ( .A(\RA2<1> ), .Y(n6) );
  INVX1 U31 ( .A(n16), .Y(n15) );
  INVX1 U32 ( .A(\RA1<2> ), .Y(n16) );
  INVX1 U33 ( .A(n8), .Y(n7) );
  INVX1 U34 ( .A(\RA2<2> ), .Y(n8) );
  INVX1 U35 ( .A(n18), .Y(n17) );
  INVX1 U36 ( .A(\RA1<3> ), .Y(n18) );
endmodule


module arm ( clk, reset, MemWrite, .Adr({\Adr<31> , \Adr<30> , \Adr<29> , 
        \Adr<28> , \Adr<27> , \Adr<26> , \Adr<25> , \Adr<24> , \Adr<23> , 
        \Adr<22> , \Adr<21> , \Adr<20> , \Adr<19> , \Adr<18> , \Adr<17> , 
        \Adr<16> , \Adr<15> , \Adr<14> , \Adr<13> , \Adr<12> , \Adr<11> , 
        \Adr<10> , \Adr<9> , \Adr<8> , \Adr<7> , \Adr<6> , \Adr<5> , \Adr<4> , 
        \Adr<3> , \Adr<2> , \Adr<1> , \Adr<0> }), .WriteData({\WriteData<31> , 
        \WriteData<30> , \WriteData<29> , \WriteData<28> , \WriteData<27> , 
        \WriteData<26> , \WriteData<25> , \WriteData<24> , \WriteData<23> , 
        \WriteData<22> , \WriteData<21> , \WriteData<20> , \WriteData<19> , 
        \WriteData<18> , \WriteData<17> , \WriteData<16> , \WriteData<15> , 
        \WriteData<14> , \WriteData<13> , \WriteData<12> , \WriteData<11> , 
        \WriteData<10> , \WriteData<9> , \WriteData<8> , \WriteData<7> , 
        \WriteData<6> , \WriteData<5> , \WriteData<4> , \WriteData<3> , 
        \WriteData<2> , \WriteData<1> , \WriteData<0> }), .ReadData({
        \ReadData<31> , \ReadData<30> , \ReadData<29> , \ReadData<28> , 
        \ReadData<27> , \ReadData<26> , \ReadData<25> , \ReadData<24> , 
        \ReadData<23> , \ReadData<22> , \ReadData<21> , \ReadData<20> , 
        \ReadData<19> , \ReadData<18> , \ReadData<17> , \ReadData<16> , 
        \ReadData<15> , \ReadData<14> , \ReadData<13> , \ReadData<12> , 
        \ReadData<11> , \ReadData<10> , \ReadData<9> , \ReadData<8> , 
        \ReadData<7> , \ReadData<6> , \ReadData<5> , \ReadData<4> , 
        \ReadData<3> , \ReadData<2> , \ReadData<1> , \ReadData<0> }) );
  input clk, reset, \ReadData<31> , \ReadData<30> , \ReadData<29> ,
         \ReadData<28> , \ReadData<27> , \ReadData<26> , \ReadData<25> ,
         \ReadData<24> , \ReadData<23> , \ReadData<22> , \ReadData<21> ,
         \ReadData<20> , \ReadData<19> , \ReadData<18> , \ReadData<17> ,
         \ReadData<16> , \ReadData<15> , \ReadData<14> , \ReadData<13> ,
         \ReadData<12> , \ReadData<11> , \ReadData<10> , \ReadData<9> ,
         \ReadData<8> , \ReadData<7> , \ReadData<6> , \ReadData<5> ,
         \ReadData<4> , \ReadData<3> , \ReadData<2> , \ReadData<1> ,
         \ReadData<0> ;
  output MemWrite, \Adr<31> , \Adr<30> , \Adr<29> , \Adr<28> , \Adr<27> ,
         \Adr<26> , \Adr<25> , \Adr<24> , \Adr<23> , \Adr<22> , \Adr<21> ,
         \Adr<20> , \Adr<19> , \Adr<18> , \Adr<17> , \Adr<16> , \Adr<15> ,
         \Adr<14> , \Adr<13> , \Adr<12> , \Adr<11> , \Adr<10> , \Adr<9> ,
         \Adr<8> , \Adr<7> , \Adr<6> , \Adr<5> , \Adr<4> , \Adr<3> , \Adr<2> ,
         \Adr<1> , \Adr<0> , \WriteData<31> , \WriteData<30> , \WriteData<29> ,
         \WriteData<28> , \WriteData<27> , \WriteData<26> , \WriteData<25> ,
         \WriteData<24> , \WriteData<23> , \WriteData<22> , \WriteData<21> ,
         \WriteData<20> , \WriteData<19> , \WriteData<18> , \WriteData<17> ,
         \WriteData<16> , \WriteData<15> , \WriteData<14> , \WriteData<13> ,
         \WriteData<12> , \WriteData<11> , \WriteData<10> , \WriteData<9> ,
         \WriteData<8> , \WriteData<7> , \WriteData<6> , \WriteData<5> ,
         \WriteData<4> , \WriteData<3> , \WriteData<2> , \WriteData<1> ,
         \WriteData<0> ;
  wire   \Instr<31> , \Instr<30> , \Instr<29> , \Instr<28> , \Instr<27> ,
         \Instr<26> , \Instr<25> , \Instr<24> , \Instr<23> , \Instr<22> ,
         \Instr<21> , \Instr<20> , \Instr<19> , \Instr<18> , \Instr<17> ,
         \Instr<16> , \Instr<15> , \Instr<14> , \Instr<13> , \Instr<12> ,
         \ALUFlags<3> , \ALUFlags<2> , \ALUFlags<1> , \ALUFlags<0> , PCWrite,
         RegWrite, IRWrite, AdrSrc, \RegSrc<1> , \RegSrc<0> , \ALUSrcA<1> ,
         \ALUSrcA<0> , \ALUSrcB<1> , \ALUSrcB<0> , \ResultSrc<1> ,
         \ResultSrc<0> , \ImmSrc<1> , \ImmSrc<0> , \ALUControl<1> ,
         \ALUControl<0> , n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12,
         n13, n14, n15;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11;

  controller c ( .clk(clk), .reset(reset), .Instr({\Instr<31> , \Instr<30> , 
        \Instr<29> , \Instr<28> , \Instr<27> , \Instr<26> , \Instr<25> , 
        \Instr<24> , \Instr<23> , \Instr<22> , \Instr<21> , \Instr<20> , 
        \Instr<19> , \Instr<18> , \Instr<17> , \Instr<16> , \Instr<15> , 
        \Instr<14> , \Instr<13> , \Instr<12> }), .ALUFlags({\ALUFlags<3> , 
        \ALUFlags<2> , \ALUFlags<1> , \ALUFlags<0> }), .PCWrite(PCWrite), 
        .MemWrite(MemWrite), .RegWrite(RegWrite), .IRWrite(IRWrite), .AdrSrc(
        AdrSrc), .RegSrc({\RegSrc<1> , \RegSrc<0> }), .ALUSrcA({\ALUSrcA<1> , 
        \ALUSrcA<0> }), .ALUSrcB({\ALUSrcB<1> , \ALUSrcB<0> }), .ResultSrc({
        \ResultSrc<1> , \ResultSrc<0> }), .ImmSrc({\ImmSrc<1> , \ImmSrc<0> }), 
        .ALUControl({\ALUControl<1> , \ALUControl<0> }) );
  datapath dp ( .clk(clk), .reset(reset), .Adr({\Adr<31> , \Adr<30> , 
        \Adr<29> , \Adr<28> , \Adr<27> , \Adr<26> , \Adr<25> , \Adr<24> , 
        \Adr<23> , \Adr<22> , \Adr<21> , \Adr<20> , \Adr<19> , \Adr<18> , 
        \Adr<17> , \Adr<16> , \Adr<15> , \Adr<14> , \Adr<13> , \Adr<12> , 
        \Adr<11> , \Adr<10> , \Adr<9> , \Adr<8> , \Adr<7> , \Adr<6> , \Adr<5> , 
        \Adr<4> , \Adr<3> , \Adr<2> , \Adr<1> , \Adr<0> }), .WriteData({
        \WriteData<31> , \WriteData<30> , \WriteData<29> , \WriteData<28> , 
        \WriteData<27> , \WriteData<26> , \WriteData<25> , \WriteData<24> , 
        \WriteData<23> , \WriteData<22> , \WriteData<21> , \WriteData<20> , 
        \WriteData<19> , \WriteData<18> , \WriteData<17> , \WriteData<16> , 
        \WriteData<15> , \WriteData<14> , \WriteData<13> , \WriteData<12> , 
        \WriteData<11> , \WriteData<10> , \WriteData<9> , \WriteData<8> , 
        \WriteData<7> , \WriteData<6> , \WriteData<5> , \WriteData<4> , 
        \WriteData<3> , \WriteData<2> , \WriteData<1> , \WriteData<0> }), 
        .ReadData({\ReadData<31> , \ReadData<30> , \ReadData<29> , 
        \ReadData<28> , \ReadData<27> , \ReadData<26> , \ReadData<25> , 
        \ReadData<24> , \ReadData<23> , \ReadData<22> , \ReadData<21> , 
        \ReadData<20> , \ReadData<19> , \ReadData<18> , \ReadData<17> , 
        \ReadData<16> , \ReadData<15> , \ReadData<14> , \ReadData<13> , 
        \ReadData<12> , \ReadData<11> , \ReadData<10> , \ReadData<9> , 
        \ReadData<8> , \ReadData<7> , \ReadData<6> , \ReadData<5> , 
        \ReadData<4> , \ReadData<3> , \ReadData<2> , \ReadData<1> , 
        \ReadData<0> }), .Instr({\Instr<31> , \Instr<30> , \Instr<29> , 
        \Instr<28> , \Instr<27> , \Instr<26> , \Instr<25> , \Instr<24> , 
        \Instr<23> , \Instr<22> , \Instr<21> , \Instr<20> , \Instr<19> , 
        \Instr<18> , \Instr<17> , \Instr<16> , \Instr<15> , \Instr<14> , 
        \Instr<13> , \Instr<12> , SYNOPSYS_UNCONNECTED__0, 
        SYNOPSYS_UNCONNECTED__1, SYNOPSYS_UNCONNECTED__2, 
        SYNOPSYS_UNCONNECTED__3, SYNOPSYS_UNCONNECTED__4, 
        SYNOPSYS_UNCONNECTED__5, SYNOPSYS_UNCONNECTED__6, 
        SYNOPSYS_UNCONNECTED__7, SYNOPSYS_UNCONNECTED__8, 
        SYNOPSYS_UNCONNECTED__9, SYNOPSYS_UNCONNECTED__10, 
        SYNOPSYS_UNCONNECTED__11}), .ALUFlags({\ALUFlags<3> , \ALUFlags<2> , 
        \ALUFlags<1> , \ALUFlags<0> }), .PCWrite(n14), .RegWrite(RegWrite), 
        .IRWrite(n12), .AdrSrc(n10), .RegSrc({\RegSrc<1> , \RegSrc<0> }), 
        .ALUSrcA({n8, n1}), .ALUSrcB({n6, \ALUSrcB<0> }), .ResultSrc({n4, 
        \ResultSrc<0> }), .ImmSrc({\ImmSrc<1> , \ImmSrc<0> }), .ALUControl({n2, 
        \ALUControl<0> }) );
  CLKINVX8 U1 ( .A(n9), .Y(n8) );
  INVX4 U2 ( .A(n7), .Y(n6) );
  CLKINVX4 U3 ( .A(\ALUSrcB<1> ), .Y(n7) );
  BUFX3 U4 ( .A(\ALUSrcA<0> ), .Y(n1) );
  INVX1 U5 ( .A(\ALUSrcA<1> ), .Y(n9) );
  INVX1 U6 ( .A(n5), .Y(n4) );
  INVX1 U7 ( .A(\ResultSrc<1> ), .Y(n5) );
  INVX1 U8 ( .A(n13), .Y(n12) );
  INVX1 U9 ( .A(IRWrite), .Y(n13) );
  INVX1 U10 ( .A(n11), .Y(n10) );
  INVX1 U11 ( .A(n15), .Y(n14) );
  INVX1 U12 ( .A(PCWrite), .Y(n15) );
  INVX1 U13 ( .A(n3), .Y(n2) );
  INVX1 U14 ( .A(\ALUControl<1> ), .Y(n3) );
  INVX1 U15 ( .A(AdrSrc), .Y(n11) );
endmodule

