
module mainfsm ( clk, reset, .Op({\Op<1> , \Op<0> }), .Funct({\Funct<5> , 
        \Funct<4> , \Funct<3> , \Funct<2> , \Funct<1> , \Funct<0> }), IRWrite, 
        AdrSrc, .ALUSrcA({\ALUSrcA<1> , \ALUSrcA<0> }), .ALUSrcB({\ALUSrcB<1> , 
        \ALUSrcB<0> }), .ResultSrc({\ResultSrc<1> , \ResultSrc<0> }), NextPC, 
        RegW, MemW, Branch, ALUOp );
  input clk, reset, \Op<1> , \Op<0> , \Funct<5> , \Funct<4> , \Funct<3> ,
         \Funct<2> , \Funct<1> , \Funct<0> ;
  output IRWrite, AdrSrc, \ALUSrcA<1> , \ALUSrcA<0> , \ALUSrcB<1> ,
         \ALUSrcB<0> , \ResultSrc<1> , \ResultSrc<0> , NextPC, RegW, MemW,
         Branch, ALUOp;
  wire   \state<3> , \state<2> , \state<1> , \state<0> , \nextstate<3> ,
         \nextstate<2> , \nextstate<1> , \nextstate<0> , n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n20, n87, n88, n89, n90, n91, n92, n93;

  DFFRHQX1 \state_reg<2>  ( .D(\nextstate<2> ), .CK(clk), .RN(n93), .Q(
        \state<2> ) );
  DFFRHQX1 \state_reg<3>  ( .D(\nextstate<3> ), .CK(clk), .RN(n93), .Q(
        \state<3> ) );
  DFFRHQX2 \state_reg<0>  ( .D(\nextstate<0> ), .CK(clk), .RN(n93), .Q(
        \state<0> ) );
  DFFRHQX2 \state_reg<1>  ( .D(\nextstate<1> ), .CK(clk), .RN(n93), .Q(
        \state<1> ) );
  NOR2X1 U3 ( .A(n89), .B(n90), .Y(\ALUSrcA<1> ) );
  BUFX3 U4 ( .A(\ALUSrcA<0> ), .Y(\ALUSrcB<1> ) );
  NAND2BX1 U5 ( .AN(\ALUSrcA<1> ), .B(n87), .Y(\ResultSrc<1> ) );
  NAND2X1 U6 ( .A(n88), .B(n89), .Y(n14) );
  INVX1 U7 ( .A(\ALUSrcA<0> ), .Y(n87) );
  INVX1 U8 ( .A(n11), .Y(ALUOp) );
  BUFX3 U9 ( .A(IRWrite), .Y(NextPC) );
  INVX1 U10 ( .A(\state<2> ), .Y(n88) );
  NOR2X1 U11 ( .A(n14), .B(\state<1> ), .Y(\ALUSrcA<0> ) );
  CLKINVX3 U12 ( .A(\state<0> ), .Y(n90) );
  INVX1 U13 ( .A(\state<3> ), .Y(n89) );
  OAI21XL U14 ( .A0(n90), .A1(n11), .B0(n20), .Y(\ALUSrcB<0> ) );
  AOI31X1 U15 ( .A0(n90), .A1(n88), .A2(\state<1> ), .B0(\ALUSrcA<1> ), .Y(n20) );
  NAND2X1 U16 ( .A(\state<2> ), .B(\state<1> ), .Y(n11) );
  NOR3X1 U17 ( .A(n90), .B(\state<1> ), .C(n88), .Y(MemW) );
  INVX1 U18 ( .A(n19), .Y(AdrSrc) );
  AOI31X1 U19 ( .A0(\state<1> ), .A1(n88), .A2(\state<0> ), .B0(MemW), .Y(n19)
         );
  NOR3X1 U20 ( .A(\state<0> ), .B(\state<1> ), .C(n88), .Y(\ResultSrc<0> ) );
  NOR2X1 U21 ( .A(n87), .B(\state<0> ), .Y(IRWrite) );
  INVX1 U22 ( .A(n18), .Y(RegW) );
  AOI21X1 U23 ( .A0(n90), .A1(\state<3> ), .B0(\ResultSrc<0> ), .Y(n18) );
  OAI21XL U24 ( .A0(n90), .A1(n15), .B0(n16), .Y(\nextstate<1> ) );
  NAND4BXL U25 ( .AN(n14), .B(\Funct<0> ), .C(\state<1> ), .D(n90), .Y(n16) );
  OAI21XL U26 ( .A0(\Op<0> ), .A1(n92), .B0(\ALUSrcA<0> ), .Y(n15) );
  INVX1 U27 ( .A(\Op<1> ), .Y(n92) );
  OAI22X1 U28 ( .A0(\state<0> ), .A1(n14), .B0(n87), .B1(n17), .Y(
        \nextstate<0> ) );
  OAI21XL U29 ( .A0(\Funct<5> ), .A1(\Op<1> ), .B0(n91), .Y(n17) );
  INVX1 U30 ( .A(\Op<0> ), .Y(n91) );
  AOI21X1 U31 ( .A0(n12), .A1(n13), .B0(n14), .Y(\nextstate<2> ) );
  NAND3X1 U32 ( .A(n91), .B(n92), .C(\state<0> ), .Y(n13) );
  OAI2BB1X1 U33 ( .A0N(n90), .A1N(\Funct<0> ), .B0(\state<1> ), .Y(n12) );
  OAI32X1 U34 ( .A0(n90), .A1(n87), .A2(n92), .B0(\state<3> ), .B1(n11), .Y(
        \nextstate<3> ) );
  INVX1 U35 ( .A(reset), .Y(n93) );
  BUFX3 U36 ( .A(\ALUSrcA<1> ), .Y(Branch) );
endmodule


module decode ( clk, reset, .Op({\Op<1> , \Op<0> }), .Funct({\Funct<5> , 
        \Funct<4> , \Funct<3> , \Funct<2> , \Funct<1> , \Funct<0> }), .Rd({
        \Rd<3> , \Rd<2> , \Rd<1> , \Rd<0> }), .FlagW({\FlagW<1> , \FlagW<0> }), 
        PCS, NextPC, RegW, MemW, IRWrite, AdrSrc, .ResultSrc({\ResultSrc<1> , 
        \ResultSrc<0> }), .ALUSrcA({\ALUSrcA<1> , \ALUSrcA<0> }), .ALUSrcB({
        \ALUSrcB<1> , \ALUSrcB<0> }), .ImmSrc({\ImmSrc<1> , \ImmSrc<0> }), 
    .RegSrc({\RegSrc<1> , \RegSrc<0> }), .ALUControl({\ALUControl<1> , 
        \ALUControl<0> }) );
  input clk, reset, \Op<1> , \Op<0> , \Funct<5> , \Funct<4> , \Funct<3> ,
         \Funct<2> , \Funct<1> , \Funct<0> , \Rd<3> , \Rd<2> , \Rd<1> ,
         \Rd<0> ;
  output \FlagW<1> , \FlagW<0> , PCS, NextPC, RegW, MemW, IRWrite, AdrSrc,
         \ResultSrc<1> , \ResultSrc<0> , \ALUSrcA<1> , \ALUSrcA<0> ,
         \ALUSrcB<1> , \ALUSrcB<0> , \ImmSrc<1> , \ImmSrc<0> , \RegSrc<1> ,
         \RegSrc<0> , \ALUControl<1> , \ALUControl<0> ;
  wire   Branch, ALUOp, n153, n151, n152, n150, n149, n4, n5, n6, n7, n139,
         n141, n143, n145, n147, n148;
  wire   SYNOPSYS_UNCONNECTED__0;

  mainfsm fsm ( .clk(clk), .reset(reset), .Op({\Op<1> , \Op<0> }), .Funct({
        \Funct<5> , \Funct<4> , \Funct<3> , \Funct<2> , \Funct<1> , \Funct<0> }), .IRWrite(n149), .AdrSrc(n150), .ALUSrcA({n152, n153}), .ALUSrcB({
        SYNOPSYS_UNCONNECTED__0, \ALUSrcB<0> }), .ResultSrc({n151, 
        \ResultSrc<0> }), .NextPC(NextPC), .RegW(RegW), .MemW(MemW), .Branch(
        Branch), .ALUOp(ALUOp) );
  BUFX3 U3 ( .A(\ALUSrcA<0> ), .Y(\ALUSrcB<1> ) );
  INVX1 U4 ( .A(n141), .Y(\ALUSrcA<0> ) );
  INVX1 U5 ( .A(n153), .Y(n141) );
  INVX1 U6 ( .A(n143), .Y(\ALUSrcA<1> ) );
  INVX1 U7 ( .A(n152), .Y(n143) );
  INVX1 U8 ( .A(ALUOp), .Y(n148) );
  INVX1 U9 ( .A(n139), .Y(\ResultSrc<1> ) );
  INVX1 U10 ( .A(n151), .Y(n139) );
  INVX1 U11 ( .A(n145), .Y(AdrSrc) );
  INVX1 U12 ( .A(n147), .Y(IRWrite) );
  INVX1 U13 ( .A(n149), .Y(n147) );
  INVX1 U14 ( .A(n6), .Y(\FlagW<1> ) );
  AOI2BB1X1 U15 ( .A0N(\Funct<4> ), .A1N(n7), .B0(n148), .Y(\ALUControl<1> )
         );
  NOR2X1 U16 ( .A(\Funct<3> ), .B(\Funct<2> ), .Y(n7) );
  AOI2BB1X1 U17 ( .A0N(\Funct<4> ), .A1N(\Funct<2> ), .B0(n148), .Y(
        \ALUControl<0> ) );
  INVX1 U18 ( .A(n150), .Y(n145) );
  INVX1 U19 ( .A(n4), .Y(PCS) );
  AOI31X1 U20 ( .A0(RegW), .A1(\Rd<3> ), .A2(n5), .B0(Branch), .Y(n4) );
  NOR3X1 U21 ( .A(n6), .B(\Funct<4> ), .C(n7), .Y(\FlagW<0> ) );
  AND3X2 U22 ( .A(\Rd<1> ), .B(\Rd<0> ), .C(\Rd<2> ), .Y(n5) );
  NAND2X1 U23 ( .A(\Funct<0> ), .B(ALUOp), .Y(n6) );
  BUFX3 U24 ( .A(\Op<1> ), .Y(\ImmSrc<1> ) );
  BUFX3 U25 ( .A(\Op<1> ), .Y(\RegSrc<0> ) );
  BUFX3 U26 ( .A(\Op<0> ), .Y(\ImmSrc<0> ) );
  BUFX3 U27 ( .A(\Op<0> ), .Y(\RegSrc<1> ) );
endmodule


module flopenr_WIDTH2_0 ( clk, reset, en, .d({\d<1> , \d<0> }), .q({\q<1> , 
        \q<0> }) );
  input clk, reset, en, \d<1> , \d<0> ;
  output \q<1> , \q<0> ;
  wire   n5, n6, n33, n34, n35, n36;

  DFFRHQX1 \q_reg<1>  ( .D(n33), .CK(clk), .RN(n36), .Q(\q<1> ) );
  DFFRHQX1 \q_reg<0>  ( .D(n34), .CK(clk), .RN(n36), .Q(\q<0> ) );
  INVX1 U2 ( .A(en), .Y(n35) );
  INVX1 U3 ( .A(n5), .Y(n33) );
  AOI22X1 U4 ( .A0(en), .A1(\d<1> ), .B0(\q<1> ), .B1(n35), .Y(n5) );
  INVX1 U5 ( .A(n6), .Y(n34) );
  AOI22X1 U6 ( .A0(\d<0> ), .A1(en), .B0(\q<0> ), .B1(n35), .Y(n6) );
  INVX1 U7 ( .A(reset), .Y(n36) );
endmodule


module flopenr_WIDTH2_1 ( clk, reset, en, .d({\d<1> , \d<0> }), .q({\q<1> , 
        \q<0> }) );
  input clk, reset, en, \d<1> , \d<0> ;
  output \q<1> , \q<0> ;
  wire   n5, n6, n35, n36, n37, n38;

  DFFRHQX1 \q_reg<1>  ( .D(n35), .CK(clk), .RN(n38), .Q(\q<1> ) );
  DFFRHQX1 \q_reg<0>  ( .D(n36), .CK(clk), .RN(n38), .Q(\q<0> ) );
  INVX1 U2 ( .A(en), .Y(n37) );
  INVX1 U3 ( .A(n6), .Y(n36) );
  AOI22X1 U4 ( .A0(\d<0> ), .A1(en), .B0(\q<0> ), .B1(n37), .Y(n6) );
  INVX1 U5 ( .A(n5), .Y(n35) );
  AOI22X1 U6 ( .A0(en), .A1(\d<1> ), .B0(\q<1> ), .B1(n37), .Y(n5) );
  INVX1 U7 ( .A(reset), .Y(n38) );
endmodule


module condcheck ( .Cond({\Cond<3> , \Cond<2> , \Cond<1> , \Cond<0> }), 
    .Flags({\Flags<3> , \Flags<2> , \Flags<1> , \Flags<0> }), CondEx );
  input \Cond<3> , \Cond<2> , \Cond<1> , \Cond<0> , \Flags<3> , \Flags<2> ,
         \Flags<1> , \Flags<0> ;
  output CondEx;
  wire   n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19,
         n40, n41, n42, n43;

  OAI21XL U2 ( .A0(n5), .A1(n41), .B0(n6), .Y(CondEx) );
  AOI222X1 U3 ( .A0(\Cond<0> ), .A1(n13), .B0(n14), .B1(n15), .C0(\Cond<1> ), 
        .C1(n16), .Y(n5) );
  AOI32X1 U4 ( .A0(\Cond<1> ), .A1(n7), .A2(\Cond<2> ), .B0(n8), .B1(n41), .Y(
        n6) );
  NOR2X1 U5 ( .A(\Flags<2> ), .B(\Cond<0> ), .Y(n14) );
  XNOR2X1 U6 ( .A(n40), .B(\Cond<0> ), .Y(n12) );
  XOR2X1 U7 ( .A(\Flags<2> ), .B(\Cond<0> ), .Y(n11) );
  OAI32X1 U8 ( .A0(n42), .A1(\Cond<1> ), .A2(n9), .B0(\Cond<2> ), .B1(n10), 
        .Y(n8) );
  XNOR2X1 U9 ( .A(\Flags<3> ), .B(\Cond<0> ), .Y(n9) );
  AOI22X1 U10 ( .A0(n11), .A1(n43), .B0(\Cond<1> ), .B1(n12), .Y(n10) );
  INVX1 U11 ( .A(\Cond<1> ), .Y(n43) );
  XOR2X1 U12 ( .A(\Flags<0> ), .B(\Flags<3> ), .Y(n17) );
  INVX1 U13 ( .A(\Cond<2> ), .Y(n42) );
  OAI21XL U14 ( .A0(\Cond<0> ), .A1(n17), .B0(n42), .Y(n16) );
  OAI21XL U15 ( .A0(\Cond<1> ), .A1(n18), .B0(n19), .Y(n13) );
  AOI21X1 U16 ( .A0(n42), .A1(n40), .B0(\Flags<2> ), .Y(n18) );
  OAI21XL U17 ( .A0(\Cond<1> ), .A1(\Cond<2> ), .B0(n17), .Y(n19) );
  INVX1 U18 ( .A(\Flags<1> ), .Y(n40) );
  XOR2X1 U19 ( .A(\Flags<0> ), .B(\Cond<0> ), .Y(n7) );
  OAI32X1 U20 ( .A0(n40), .A1(\Cond<2> ), .A2(\Cond<1> ), .B0(n42), .B1(n17), 
        .Y(n15) );
  INVX1 U21 ( .A(\Cond<3> ), .Y(n41) );
endmodule


module flopr_WIDTH1 ( clk, reset, .d(\d<0> ), .q(\q<0> ) );
  input clk, reset, \d<0> ;
  output \q<0> ;
  wire   n7;

  DFFRHQX1 \q_reg<0>  ( .D(\d<0> ), .CK(clk), .RN(n7), .Q(\q<0> ) );
  INVXL U3 ( .A(reset), .Y(n7) );
endmodule


module condlogic ( clk, reset, .Cond({\Cond<3> , \Cond<2> , \Cond<1> , 
        \Cond<0> }), .ALUFlags({\ALUFlags<3> , \ALUFlags<2> , \ALUFlags<1> , 
        \ALUFlags<0> }), .FlagW({\FlagW<1> , \FlagW<0> }), PCS, NextPC, RegW, 
        MemW, PCWrite, RegWrite, MemWrite );
  input clk, reset, \Cond<3> , \Cond<2> , \Cond<1> , \Cond<0> , \ALUFlags<3> ,
         \ALUFlags<2> , \ALUFlags<1> , \ALUFlags<0> , \FlagW<1> , \FlagW<0> ,
         PCS, NextPC, RegW, MemW;
  output PCWrite, RegWrite, MemWrite;
  wire   \FlagWrite<1> , \FlagWrite<0> , \Flags<3> , \Flags<2> , \Flags<1> ,
         \Flags<0> , CondEx, CondExDelayed, n2;

  flopenr_WIDTH2_0 flagreg1 ( .clk(clk), .reset(reset), .en(\FlagWrite<1> ), 
        .d({\ALUFlags<3> , \ALUFlags<2> }), .q({\Flags<3> , \Flags<2> }) );
  flopenr_WIDTH2_1 flagreg0 ( .clk(clk), .reset(reset), .en(\FlagWrite<0> ), 
        .d({\ALUFlags<1> , \ALUFlags<0> }), .q({\Flags<1> , \Flags<0> }) );
  condcheck cc ( .Cond({\Cond<3> , \Cond<2> , \Cond<1> , \Cond<0> }), .Flags({
        \Flags<3> , \Flags<2> , \Flags<1> , \Flags<0> }), .CondEx(CondEx) );
  flopr_WIDTH1 condreg ( .clk(clk), .reset(reset), .d(CondEx), .q(
        CondExDelayed) );
  AND2X2 U1 ( .A(\FlagW<1> ), .B(CondEx), .Y(\FlagWrite<1> ) );
  INVX1 U2 ( .A(n2), .Y(PCWrite) );
  AOI21X1 U3 ( .A0(PCS), .A1(CondExDelayed), .B0(NextPC), .Y(n2) );
  AND2X2 U4 ( .A(RegW), .B(CondExDelayed), .Y(RegWrite) );
  AND2X2 U5 ( .A(\FlagW<0> ), .B(CondEx), .Y(\FlagWrite<0> ) );
  AND2X2 U6 ( .A(MemW), .B(CondExDelayed), .Y(MemWrite) );
endmodule


module controller ( clk, reset, .Instr({\Instr<31> , \Instr<30> , \Instr<29> , 
        \Instr<28> , \Instr<27> , \Instr<26> , \Instr<25> , \Instr<24> , 
        \Instr<23> , \Instr<22> , \Instr<21> , \Instr<20> , \Instr<19> , 
        \Instr<18> , \Instr<17> , \Instr<16> , \Instr<15> , \Instr<14> , 
        \Instr<13> , \Instr<12> }), .ALUFlags({\ALUFlags<3> , \ALUFlags<2> , 
        \ALUFlags<1> , \ALUFlags<0> }), PCWrite, MemWrite, RegWrite, IRWrite, 
        AdrSrc, .RegSrc({\RegSrc<1> , \RegSrc<0> }), .ALUSrcA({\ALUSrcA<1> , 
        \ALUSrcA<0> }), .ALUSrcB({\ALUSrcB<1> , \ALUSrcB<0> }), .ResultSrc({
        \ResultSrc<1> , \ResultSrc<0> }), .ImmSrc({\ImmSrc<1> , \ImmSrc<0> }), 
    .ALUControl({\ALUControl<1> , \ALUControl<0> }) );
  input clk, reset, \Instr<31> , \Instr<30> , \Instr<29> , \Instr<28> ,
         \Instr<27> , \Instr<26> , \Instr<25> , \Instr<24> , \Instr<23> ,
         \Instr<22> , \Instr<21> , \Instr<20> , \Instr<19> , \Instr<18> ,
         \Instr<17> , \Instr<16> , \Instr<15> , \Instr<14> , \Instr<13> ,
         \Instr<12> , \ALUFlags<3> , \ALUFlags<2> , \ALUFlags<1> ,
         \ALUFlags<0> ;
  output PCWrite, MemWrite, RegWrite, IRWrite, AdrSrc, \RegSrc<1> ,
         \RegSrc<0> , \ALUSrcA<1> , \ALUSrcA<0> , \ALUSrcB<1> , \ALUSrcB<0> ,
         \ResultSrc<1> , \ResultSrc<0> , \ImmSrc<1> , \ImmSrc<0> ,
         \ALUControl<1> , \ALUControl<0> ;
  wire   \FlagW<1> , \FlagW<0> , PCS, RegW, MemW, n153, n152, n151, n150, n149,
         n148, n147, n134, n136, n138, n140, n142, n144, n146;

  decode dec ( .clk(clk), .reset(reset), .Op({\Instr<27> , \Instr<26> }), 
        .Funct({\Instr<25> , \Instr<24> , \Instr<23> , \Instr<22> , 
        \Instr<21> , \Instr<20> }), .Rd({\Instr<15> , \Instr<14> , \Instr<13> , 
        \Instr<12> }), .FlagW({\FlagW<1> , \FlagW<0> }), .PCS(PCS), .RegW(RegW), .MemW(MemW), .IRWrite(n148), .AdrSrc(n149), .ResultSrc({n152, \ResultSrc<0> }), .ALUSrcA({n150, n151}), .ALUSrcB({\ALUSrcB<1> , \ALUSrcB<0> }), .ImmSrc({
        \ImmSrc<1> , \ImmSrc<0> }), .RegSrc({\RegSrc<1> , \RegSrc<0> }), 
        .ALUControl({n153, \ALUControl<0> }) );
  condlogic cl ( .clk(clk), .reset(reset), .Cond({\Instr<31> , \Instr<30> , 
        \Instr<29> , \Instr<28> }), .ALUFlags({\ALUFlags<3> , \ALUFlags<2> , 
        \ALUFlags<1> , \ALUFlags<0> }), .FlagW({\FlagW<1> , \FlagW<0> }), 
        .PCS(PCS), .NextPC(IRWrite), .RegW(RegW), .MemW(MemW), .PCWrite(n147), 
        .RegWrite(RegWrite), .MemWrite(MemWrite) );
  INVX1 U1 ( .A(n138), .Y(\ALUSrcA<0> ) );
  INVX1 U2 ( .A(n151), .Y(n138) );
  INVX1 U3 ( .A(n140), .Y(\ALUSrcA<1> ) );
  INVX1 U4 ( .A(n150), .Y(n140) );
  INVX1 U5 ( .A(n136), .Y(\ResultSrc<1> ) );
  INVX1 U6 ( .A(n152), .Y(n136) );
  INVX1 U7 ( .A(n134), .Y(\ALUControl<1> ) );
  INVX1 U8 ( .A(n153), .Y(n134) );
  INVX1 U9 ( .A(n142), .Y(AdrSrc) );
  INVX1 U10 ( .A(n149), .Y(n142) );
  INVX1 U11 ( .A(n144), .Y(IRWrite) );
  INVX1 U12 ( .A(n148), .Y(n144) );
  INVX1 U13 ( .A(n146), .Y(PCWrite) );
  INVX1 U14 ( .A(n147), .Y(n146) );
endmodule


module flopenr_WIDTH32_0 ( clk, reset, en, .d({\d<31> , \d<30> , \d<29> , 
        \d<28> , \d<27> , \d<26> , \d<25> , \d<24> , \d<23> , \d<22> , \d<21> , 
        \d<20> , \d<19> , \d<18> , \d<17> , \d<16> , \d<15> , \d<14> , \d<13> , 
        \d<12> , \d<11> , \d<10> , \d<9> , \d<8> , \d<7> , \d<6> , \d<5> , 
        \d<4> , \d<3> , \d<2> , \d<1> , \d<0> }), .q({\q<31> , \q<30> , 
        \q<29> , \q<28> , \q<27> , \q<26> , \q<25> , \q<24> , \q<23> , \q<22> , 
        \q<21> , \q<20> , \q<19> , \q<18> , \q<17> , \q<16> , \q<15> , \q<14> , 
        \q<13> , \q<12> , \q<11> , \q<10> , \q<9> , \q<8> , \q<7> , \q<6> , 
        \q<5> , \q<4> , \q<3> , \q<2> , \q<1> , \q<0> }) );
  input clk, reset, en, \d<31> , \d<30> , \d<29> , \d<28> , \d<27> , \d<26> ,
         \d<25> , \d<24> , \d<23> , \d<22> , \d<21> , \d<20> , \d<19> ,
         \d<18> , \d<17> , \d<16> , \d<15> , \d<14> , \d<13> , \d<12> ,
         \d<11> , \d<10> , \d<9> , \d<8> , \d<7> , \d<6> , \d<5> , \d<4> ,
         \d<3> , \d<2> , \d<1> , \d<0> ;
  output \q<31> , \q<30> , \q<29> , \q<28> , \q<27> , \q<26> , \q<25> ,
         \q<24> , \q<23> , \q<22> , \q<21> , \q<20> , \q<19> , \q<18> ,
         \q<17> , \q<16> , \q<15> , \q<14> , \q<13> , \q<12> , \q<11> ,
         \q<10> , \q<9> , \q<8> , \q<7> , \q<6> , \q<5> , \q<4> , \q<3> ,
         \q<2> , \q<1> , \q<0> ;
  wire   n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62,
         n63, n64, n65, n66, n301, n302, n303, n304, n305, n306, n307, n308,
         n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319,
         n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330,
         n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341,
         n342, n343, n344, n345;

  DFFRHQX1 \q_reg<31>  ( .D(n313), .CK(clk), .RN(n301), .Q(\q<31> ) );
  DFFRHQX1 \q_reg<30>  ( .D(n314), .CK(clk), .RN(n302), .Q(\q<30> ) );
  DFFRHQX1 \q_reg<29>  ( .D(n315), .CK(clk), .RN(n301), .Q(\q<29> ) );
  DFFRHQX1 \q_reg<28>  ( .D(n316), .CK(clk), .RN(n302), .Q(\q<28> ) );
  DFFRHQX1 \q_reg<27>  ( .D(n317), .CK(clk), .RN(n301), .Q(\q<27> ) );
  DFFRHQX1 \q_reg<26>  ( .D(n318), .CK(clk), .RN(n302), .Q(\q<26> ) );
  DFFRHQX1 \q_reg<25>  ( .D(n319), .CK(clk), .RN(n345), .Q(\q<25> ) );
  DFFRHQX1 \q_reg<24>  ( .D(n320), .CK(clk), .RN(n345), .Q(\q<24> ) );
  DFFRHQX1 \q_reg<23>  ( .D(n321), .CK(clk), .RN(n302), .Q(\q<23> ) );
  DFFRHQX1 \q_reg<22>  ( .D(n322), .CK(clk), .RN(n302), .Q(\q<22> ) );
  DFFRHQX1 \q_reg<21>  ( .D(n323), .CK(clk), .RN(n302), .Q(\q<21> ) );
  DFFRHQX1 \q_reg<20>  ( .D(n324), .CK(clk), .RN(n302), .Q(\q<20> ) );
  DFFRHQX1 \q_reg<19>  ( .D(n325), .CK(clk), .RN(n302), .Q(\q<19> ) );
  DFFRHQX1 \q_reg<18>  ( .D(n326), .CK(clk), .RN(n302), .Q(\q<18> ) );
  DFFRHQX1 \q_reg<17>  ( .D(n327), .CK(clk), .RN(n302), .Q(\q<17> ) );
  DFFRHQX1 \q_reg<16>  ( .D(n328), .CK(clk), .RN(n302), .Q(\q<16> ) );
  DFFRHQX1 \q_reg<15>  ( .D(n329), .CK(clk), .RN(n302), .Q(\q<15> ) );
  DFFRHQX1 \q_reg<14>  ( .D(n330), .CK(clk), .RN(n302), .Q(\q<14> ) );
  DFFRHQX1 \q_reg<13>  ( .D(n331), .CK(clk), .RN(n302), .Q(\q<13> ) );
  DFFRHQX1 \q_reg<12>  ( .D(n332), .CK(clk), .RN(n302), .Q(\q<12> ) );
  DFFRHQX1 \q_reg<11>  ( .D(n333), .CK(clk), .RN(n301), .Q(\q<11> ) );
  DFFRHQX1 \q_reg<10>  ( .D(n334), .CK(clk), .RN(n301), .Q(\q<10> ) );
  DFFRHQX1 \q_reg<9>  ( .D(n335), .CK(clk), .RN(n301), .Q(\q<9> ) );
  DFFRHQX1 \q_reg<8>  ( .D(n336), .CK(clk), .RN(n301), .Q(\q<8> ) );
  DFFRHQX1 \q_reg<7>  ( .D(n337), .CK(clk), .RN(n301), .Q(\q<7> ) );
  DFFRHQX1 \q_reg<6>  ( .D(n338), .CK(clk), .RN(n301), .Q(\q<6> ) );
  DFFRHQX1 \q_reg<5>  ( .D(n339), .CK(clk), .RN(n301), .Q(\q<5> ) );
  DFFRHQX1 \q_reg<4>  ( .D(n340), .CK(clk), .RN(n301), .Q(\q<4> ) );
  DFFRHQX1 \q_reg<3>  ( .D(n341), .CK(clk), .RN(n301), .Q(\q<3> ) );
  DFFRHQX1 \q_reg<2>  ( .D(n342), .CK(clk), .RN(n301), .Q(\q<2> ) );
  DFFRHQX1 \q_reg<1>  ( .D(n343), .CK(clk), .RN(n301), .Q(\q<1> ) );
  DFFRHQX1 \q_reg<0>  ( .D(n344), .CK(clk), .RN(n301), .Q(\q<0> ) );
  CLKINVX3 U2 ( .A(n312), .Y(n304) );
  INVX1 U3 ( .A(n310), .Y(n309) );
  INVX1 U4 ( .A(n310), .Y(n308) );
  INVX1 U5 ( .A(n311), .Y(n307) );
  INVX1 U6 ( .A(n311), .Y(n306) );
  INVX1 U7 ( .A(n311), .Y(n305) );
  INVX1 U8 ( .A(n312), .Y(n310) );
  INVX1 U9 ( .A(n312), .Y(n311) );
  INVX1 U10 ( .A(en), .Y(n312) );
  CLKINVX3 U11 ( .A(n303), .Y(n302) );
  CLKINVX3 U12 ( .A(n303), .Y(n301) );
  INVX1 U13 ( .A(n345), .Y(n303) );
  INVX1 U14 ( .A(n35), .Y(n313) );
  AOI22X1 U15 ( .A0(n311), .A1(\d<31> ), .B0(\q<31> ), .B1(n305), .Y(n35) );
  INVX1 U16 ( .A(n38), .Y(n316) );
  AOI22X1 U17 ( .A0(\d<28> ), .A1(n310), .B0(\q<28> ), .B1(n306), .Y(n38) );
  INVX1 U18 ( .A(n37), .Y(n315) );
  AOI22X1 U19 ( .A0(\d<29> ), .A1(en), .B0(\q<29> ), .B1(n306), .Y(n37) );
  INVX1 U20 ( .A(n36), .Y(n314) );
  AOI22X1 U21 ( .A0(\d<30> ), .A1(n311), .B0(\q<30> ), .B1(n305), .Y(n36) );
  INVX1 U22 ( .A(n43), .Y(n321) );
  AOI22X1 U23 ( .A0(\d<23> ), .A1(n304), .B0(\q<23> ), .B1(n308), .Y(n43) );
  INVX1 U24 ( .A(n42), .Y(n320) );
  AOI22X1 U25 ( .A0(\d<24> ), .A1(n311), .B0(\q<24> ), .B1(n309), .Y(n42) );
  INVX1 U26 ( .A(n41), .Y(n319) );
  AOI22X1 U27 ( .A0(\d<25> ), .A1(n304), .B0(\q<25> ), .B1(n305), .Y(n41) );
  INVX1 U28 ( .A(n40), .Y(n318) );
  AOI22X1 U29 ( .A0(\d<26> ), .A1(n310), .B0(\q<26> ), .B1(n307), .Y(n40) );
  INVX1 U30 ( .A(n39), .Y(n317) );
  AOI22X1 U31 ( .A0(\d<27> ), .A1(en), .B0(\q<27> ), .B1(n307), .Y(n39) );
  INVX1 U32 ( .A(n48), .Y(n326) );
  AOI22X1 U33 ( .A0(\d<18> ), .A1(n304), .B0(\q<18> ), .B1(n308), .Y(n48) );
  INVX1 U34 ( .A(n47), .Y(n325) );
  AOI22X1 U35 ( .A0(\d<19> ), .A1(n304), .B0(\q<19> ), .B1(n309), .Y(n47) );
  INVX1 U36 ( .A(n46), .Y(n324) );
  AOI22X1 U37 ( .A0(\d<20> ), .A1(n304), .B0(\q<20> ), .B1(n308), .Y(n46) );
  INVX1 U38 ( .A(n45), .Y(n323) );
  AOI22X1 U39 ( .A0(\d<21> ), .A1(n304), .B0(\q<21> ), .B1(n308), .Y(n45) );
  INVX1 U40 ( .A(n44), .Y(n322) );
  AOI22X1 U41 ( .A0(\d<22> ), .A1(n304), .B0(\q<22> ), .B1(n306), .Y(n44) );
  INVX1 U42 ( .A(n53), .Y(n331) );
  AOI22X1 U43 ( .A0(\d<13> ), .A1(n304), .B0(\q<13> ), .B1(n307), .Y(n53) );
  INVX1 U44 ( .A(n52), .Y(n330) );
  AOI22X1 U45 ( .A0(\d<14> ), .A1(n311), .B0(\q<14> ), .B1(n312), .Y(n52) );
  INVX1 U46 ( .A(n51), .Y(n329) );
  AOI22X1 U47 ( .A0(\d<15> ), .A1(n310), .B0(\q<15> ), .B1(n308), .Y(n51) );
  INVX1 U48 ( .A(n50), .Y(n328) );
  AOI22X1 U49 ( .A0(\d<16> ), .A1(n310), .B0(\q<16> ), .B1(n308), .Y(n50) );
  INVX1 U50 ( .A(n49), .Y(n327) );
  AOI22X1 U51 ( .A0(\d<17> ), .A1(en), .B0(\q<17> ), .B1(n312), .Y(n49) );
  INVX1 U52 ( .A(n58), .Y(n336) );
  AOI22X1 U53 ( .A0(\d<8> ), .A1(n304), .B0(\q<8> ), .B1(n306), .Y(n58) );
  INVX1 U54 ( .A(n57), .Y(n335) );
  AOI22X1 U55 ( .A0(\d<9> ), .A1(n304), .B0(\q<9> ), .B1(n308), .Y(n57) );
  INVX1 U56 ( .A(n56), .Y(n334) );
  AOI22X1 U57 ( .A0(\d<10> ), .A1(n304), .B0(\q<10> ), .B1(n309), .Y(n56) );
  INVX1 U58 ( .A(n55), .Y(n333) );
  AOI22X1 U59 ( .A0(\d<11> ), .A1(n304), .B0(\q<11> ), .B1(n309), .Y(n55) );
  INVX1 U60 ( .A(n54), .Y(n332) );
  AOI22X1 U61 ( .A0(\d<12> ), .A1(en), .B0(\q<12> ), .B1(n305), .Y(n54) );
  INVX1 U62 ( .A(n64), .Y(n342) );
  AOI22X1 U63 ( .A0(\d<2> ), .A1(n304), .B0(\q<2> ), .B1(n312), .Y(n64) );
  INVX1 U64 ( .A(n63), .Y(n341) );
  AOI22X1 U65 ( .A0(\d<3> ), .A1(n304), .B0(\q<3> ), .B1(n307), .Y(n63) );
  INVX1 U66 ( .A(n62), .Y(n340) );
  AOI22X1 U67 ( .A0(\d<4> ), .A1(n304), .B0(\q<4> ), .B1(n306), .Y(n62) );
  INVX1 U68 ( .A(n61), .Y(n339) );
  AOI22X1 U69 ( .A0(\d<5> ), .A1(n304), .B0(\q<5> ), .B1(n305), .Y(n61) );
  INVX1 U70 ( .A(n60), .Y(n338) );
  AOI22X1 U71 ( .A0(\d<6> ), .A1(n304), .B0(\q<6> ), .B1(n309), .Y(n60) );
  INVX1 U72 ( .A(n59), .Y(n337) );
  AOI22X1 U73 ( .A0(\d<7> ), .A1(n304), .B0(\q<7> ), .B1(n309), .Y(n59) );
  INVX1 U74 ( .A(n66), .Y(n344) );
  AOI22X1 U75 ( .A0(\d<0> ), .A1(n304), .B0(\q<0> ), .B1(n307), .Y(n66) );
  INVX1 U76 ( .A(n65), .Y(n343) );
  AOI22X1 U77 ( .A0(\d<1> ), .A1(n304), .B0(\q<1> ), .B1(n309), .Y(n65) );
  INVXL U78 ( .A(reset), .Y(n345) );
endmodule


module flopenr_WIDTH32_1 ( clk, reset, en, .d({\d<31> , \d<30> , \d<29> , 
        \d<28> , \d<27> , \d<26> , \d<25> , \d<24> , \d<23> , \d<22> , \d<21> , 
        \d<20> , \d<19> , \d<18> , \d<17> , \d<16> , \d<15> , \d<14> , \d<13> , 
        \d<12> , \d<11> , \d<10> , \d<9> , \d<8> , \d<7> , \d<6> , \d<5> , 
        \d<4> , \d<3> , \d<2> , \d<1> , \d<0> }), .q({\q<31> , \q<30> , 
        \q<29> , \q<28> , \q<27> , \q<26> , \q<25> , \q<24> , \q<23> , \q<22> , 
        \q<21> , \q<20> , \q<19> , \q<18> , \q<17> , \q<16> , \q<15> , \q<14> , 
        \q<13> , \q<12> , \q<11> , \q<10> , \q<9> , \q<8> , \q<7> , \q<6> , 
        \q<5> , \q<4> , \q<3> , \q<2> , \q<1> , \q<0> }) );
  input clk, reset, en, \d<31> , \d<30> , \d<29> , \d<28> , \d<27> , \d<26> ,
         \d<25> , \d<24> , \d<23> , \d<22> , \d<21> , \d<20> , \d<19> ,
         \d<18> , \d<17> , \d<16> , \d<15> , \d<14> , \d<13> , \d<12> ,
         \d<11> , \d<10> , \d<9> , \d<8> , \d<7> , \d<6> , \d<5> , \d<4> ,
         \d<3> , \d<2> , \d<1> , \d<0> ;
  output \q<31> , \q<30> , \q<29> , \q<28> , \q<27> , \q<26> , \q<25> ,
         \q<24> , \q<23> , \q<22> , \q<21> , \q<20> , \q<19> , \q<18> ,
         \q<17> , \q<16> , \q<15> , \q<14> , \q<13> , \q<12> , \q<11> ,
         \q<10> , \q<9> , \q<8> , \q<7> , \q<6> , \q<5> , \q<4> , \q<3> ,
         \q<2> , \q<1> , \q<0> ;
  wire   n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62,
         n63, n64, n65, n66, n333, n334, n335, n336, n337, n338, n339, n340,
         n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351,
         n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362,
         n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373,
         n374, n375, n376, n377;

  DFFRHQX1 \q_reg<25>  ( .D(n362), .CK(clk), .RN(n334), .Q(\q<25> ) );
  DFFRHQX1 \q_reg<31>  ( .D(n369), .CK(clk), .RN(n333), .Q(\q<31> ) );
  DFFRHQX2 \q_reg<30>  ( .D(n368), .CK(clk), .RN(n333), .Q(\q<30> ) );
  DFFRHQX1 \q_reg<21>  ( .D(n358), .CK(clk), .RN(n334), .Q(\q<21> ) );
  DFFRHQX1 \q_reg<23>  ( .D(n360), .CK(clk), .RN(n333), .Q(\q<23> ) );
  DFFRHQX1 \q_reg<19>  ( .D(n355), .CK(clk), .RN(n334), .Q(\q<19> ) );
  DFFRHQX1 \q_reg<18>  ( .D(n354), .CK(clk), .RN(n377), .Q(\q<18> ) );
  DFFRHQX1 \q_reg<17>  ( .D(n353), .CK(clk), .RN(n377), .Q(\q<17> ) );
  DFFRHQX1 \q_reg<22>  ( .D(n359), .CK(clk), .RN(n334), .Q(\q<22> ) );
  DFFRHQX1 \q_reg<24>  ( .D(n361), .CK(clk), .RN(n334), .Q(\q<24> ) );
  DFFRHQX1 \q_reg<16>  ( .D(n352), .CK(clk), .RN(n334), .Q(\q<16> ) );
  DFFRHQX2 \q_reg<14>  ( .D(n350), .CK(clk), .RN(n334), .Q(\q<14> ) );
  DFFRHQX2 \q_reg<15>  ( .D(n351), .CK(clk), .RN(n334), .Q(\q<15> ) );
  DFFRHQX1 \q_reg<11>  ( .D(n347), .CK(clk), .RN(n334), .Q(\q<11> ) );
  DFFRHQX1 \q_reg<10>  ( .D(n346), .CK(clk), .RN(n334), .Q(\q<10> ) );
  DFFRHQX2 \q_reg<12>  ( .D(n348), .CK(clk), .RN(n334), .Q(\q<12> ) );
  DFFRHQX2 \q_reg<13>  ( .D(n349), .CK(clk), .RN(n334), .Q(\q<13> ) );
  DFFRHQX1 \q_reg<9>  ( .D(n376), .CK(clk), .RN(n334), .Q(\q<9> ) );
  DFFRHQX1 \q_reg<8>  ( .D(n375), .CK(clk), .RN(n334), .Q(\q<8> ) );
  DFFRHQX1 \q_reg<7>  ( .D(n374), .CK(clk), .RN(n333), .Q(\q<7> ) );
  DFFRHQX1 \q_reg<6>  ( .D(n373), .CK(clk), .RN(n333), .Q(\q<6> ) );
  DFFRHQX1 \q_reg<5>  ( .D(n372), .CK(clk), .RN(n333), .Q(\q<5> ) );
  DFFRHQX1 \q_reg<4>  ( .D(n371), .CK(clk), .RN(n333), .Q(\q<4> ) );
  DFFRHQX1 \q_reg<3>  ( .D(n370), .CK(clk), .RN(n333), .Q(\q<3> ) );
  DFFRHQX1 \q_reg<2>  ( .D(n367), .CK(clk), .RN(n333), .Q(\q<2> ) );
  DFFRHQX1 \q_reg<1>  ( .D(n356), .CK(clk), .RN(n333), .Q(\q<1> ) );
  DFFRHQX1 \q_reg<0>  ( .D(n345), .CK(clk), .RN(n333), .Q(\q<0> ) );
  DFFRHQX1 \q_reg<20>  ( .D(n357), .CK(clk), .RN(n334), .Q(\q<20> ) );
  DFFRHQX1 \q_reg<26>  ( .D(n363), .CK(clk), .RN(n333), .Q(\q<26> ) );
  DFFRHQX1 \q_reg<27>  ( .D(n364), .CK(clk), .RN(n333), .Q(\q<27> ) );
  DFFRHQX2 \q_reg<29>  ( .D(n366), .CK(clk), .RN(n333), .Q(\q<29> ) );
  DFFRHQX2 \q_reg<28>  ( .D(n365), .CK(clk), .RN(n333), .Q(\q<28> ) );
  CLKINVX3 U2 ( .A(n344), .Y(n336) );
  INVX1 U3 ( .A(n342), .Y(n341) );
  INVX1 U4 ( .A(n342), .Y(n340) );
  INVX1 U5 ( .A(n343), .Y(n339) );
  INVX1 U6 ( .A(n343), .Y(n338) );
  INVX1 U7 ( .A(n343), .Y(n337) );
  INVX1 U8 ( .A(n344), .Y(n342) );
  INVX1 U9 ( .A(n344), .Y(n343) );
  INVX1 U10 ( .A(en), .Y(n344) );
  CLKINVX3 U11 ( .A(n335), .Y(n334) );
  CLKINVX3 U12 ( .A(n335), .Y(n333) );
  INVX1 U13 ( .A(n377), .Y(n335) );
  INVX1 U14 ( .A(n35), .Y(n362) );
  AOI22X1 U15 ( .A0(n342), .A1(\d<25> ), .B0(\q<25> ), .B1(n337), .Y(n35) );
  INVX1 U16 ( .A(n66), .Y(n365) );
  AOI22X1 U17 ( .A0(\d<28> ), .A1(n336), .B0(\q<28> ), .B1(n341), .Y(n66) );
  INVX1 U18 ( .A(n65), .Y(n366) );
  AOI22X1 U19 ( .A0(\d<29> ), .A1(n336), .B0(\q<29> ), .B1(n337), .Y(n65) );
  INVX1 U20 ( .A(n48), .Y(n351) );
  AOI22X1 U21 ( .A0(\d<15> ), .A1(n336), .B0(\q<15> ), .B1(n338), .Y(n48) );
  INVX1 U22 ( .A(n47), .Y(n350) );
  AOI22X1 U23 ( .A0(\d<14> ), .A1(n336), .B0(\q<14> ), .B1(n338), .Y(n47) );
  INVX1 U24 ( .A(n52), .Y(n349) );
  AOI22X1 U25 ( .A0(\d<13> ), .A1(n336), .B0(\q<13> ), .B1(n339), .Y(n52) );
  INVX1 U26 ( .A(n51), .Y(n348) );
  AOI22X1 U27 ( .A0(\d<12> ), .A1(n336), .B0(\q<12> ), .B1(n339), .Y(n51) );
  INVX1 U28 ( .A(n37), .Y(n368) );
  AOI22X1 U29 ( .A0(\d<30> ), .A1(n336), .B0(\q<30> ), .B1(n337), .Y(n37) );
  INVX1 U30 ( .A(n63), .Y(n363) );
  AOI22X1 U31 ( .A0(\d<26> ), .A1(n336), .B0(\q<26> ), .B1(n339), .Y(n63) );
  INVX1 U32 ( .A(n64), .Y(n364) );
  AOI22X1 U33 ( .A0(\d<27> ), .A1(n336), .B0(\q<27> ), .B1(n338), .Y(n64) );
  INVX1 U34 ( .A(n45), .Y(n357) );
  AOI22X1 U35 ( .A0(\d<20> ), .A1(n343), .B0(\q<20> ), .B1(n340), .Y(n45) );
  INVX1 U36 ( .A(n62), .Y(n345) );
  AOI22X1 U37 ( .A0(\d<0> ), .A1(n336), .B0(\q<0> ), .B1(n341), .Y(n62) );
  INVX1 U38 ( .A(n61), .Y(n356) );
  AOI22X1 U39 ( .A0(\d<1> ), .A1(n336), .B0(\q<1> ), .B1(n340), .Y(n61) );
  INVX1 U40 ( .A(n60), .Y(n367) );
  AOI22X1 U41 ( .A0(\d<2> ), .A1(n336), .B0(\q<2> ), .B1(n337), .Y(n60) );
  INVX1 U42 ( .A(n59), .Y(n370) );
  AOI22X1 U43 ( .A0(\d<3> ), .A1(n336), .B0(\q<3> ), .B1(n339), .Y(n59) );
  INVX1 U44 ( .A(n58), .Y(n371) );
  AOI22X1 U45 ( .A0(\d<4> ), .A1(n336), .B0(\q<4> ), .B1(n341), .Y(n58) );
  INVX1 U46 ( .A(n57), .Y(n372) );
  AOI22X1 U47 ( .A0(\d<5> ), .A1(n336), .B0(\q<5> ), .B1(n341), .Y(n57) );
  INVX1 U48 ( .A(n56), .Y(n373) );
  AOI22X1 U49 ( .A0(\d<6> ), .A1(n336), .B0(\q<6> ), .B1(n340), .Y(n56) );
  INVX1 U50 ( .A(n55), .Y(n374) );
  AOI22X1 U51 ( .A0(\d<7> ), .A1(n336), .B0(\q<7> ), .B1(n340), .Y(n55) );
  INVX1 U52 ( .A(n54), .Y(n375) );
  AOI22X1 U53 ( .A0(\d<8> ), .A1(en), .B0(\q<8> ), .B1(n341), .Y(n54) );
  INVX1 U54 ( .A(n53), .Y(n376) );
  AOI22X1 U55 ( .A0(\d<9> ), .A1(en), .B0(\q<9> ), .B1(n340), .Y(n53) );
  INVX1 U56 ( .A(n50), .Y(n346) );
  AOI22X1 U57 ( .A0(\d<10> ), .A1(en), .B0(\q<10> ), .B1(n338), .Y(n50) );
  INVX1 U58 ( .A(n49), .Y(n347) );
  AOI22X1 U59 ( .A0(\d<11> ), .A1(en), .B0(\q<11> ), .B1(n339), .Y(n49) );
  INVX1 U60 ( .A(n46), .Y(n352) );
  AOI22X1 U61 ( .A0(\d<16> ), .A1(en), .B0(\q<16> ), .B1(n344), .Y(n46) );
  INVX1 U62 ( .A(n44), .Y(n361) );
  AOI22X1 U63 ( .A0(\d<24> ), .A1(n336), .B0(\q<24> ), .B1(n341), .Y(n44) );
  INVX1 U64 ( .A(n43), .Y(n359) );
  AOI22X1 U65 ( .A0(\d<22> ), .A1(n342), .B0(\q<22> ), .B1(n344), .Y(n43) );
  INVX1 U66 ( .A(n42), .Y(n353) );
  AOI22X1 U67 ( .A0(\d<17> ), .A1(n343), .B0(\q<17> ), .B1(n341), .Y(n42) );
  INVX1 U68 ( .A(n41), .Y(n354) );
  AOI22X1 U69 ( .A0(\d<18> ), .A1(n336), .B0(\q<18> ), .B1(n340), .Y(n41) );
  INVX1 U70 ( .A(n40), .Y(n355) );
  AOI22X1 U71 ( .A0(\d<19> ), .A1(n342), .B0(\q<19> ), .B1(n340), .Y(n40) );
  INVX1 U72 ( .A(n39), .Y(n360) );
  AOI22X1 U73 ( .A0(\d<23> ), .A1(n342), .B0(\q<23> ), .B1(n338), .Y(n39) );
  INVX1 U74 ( .A(n38), .Y(n358) );
  AOI22X1 U75 ( .A0(\d<21> ), .A1(n343), .B0(\q<21> ), .B1(n339), .Y(n38) );
  INVX1 U76 ( .A(n36), .Y(n369) );
  AOI22X1 U77 ( .A0(\d<31> ), .A1(n336), .B0(\q<31> ), .B1(n337), .Y(n36) );
  INVXL U78 ( .A(reset), .Y(n377) );
endmodule


module flopr_WIDTH32_0 ( clk, reset, .d({\d<31> , \d<30> , \d<29> , \d<28> , 
        \d<27> , \d<26> , \d<25> , \d<24> , \d<23> , \d<22> , \d<21> , \d<20> , 
        \d<19> , \d<18> , \d<17> , \d<16> , \d<15> , \d<14> , \d<13> , \d<12> , 
        \d<11> , \d<10> , \d<9> , \d<8> , \d<7> , \d<6> , \d<5> , \d<4> , 
        \d<3> , \d<2> , \d<1> , \d<0> }), .q({\q<31> , \q<30> , \q<29> , 
        \q<28> , \q<27> , \q<26> , \q<25> , \q<24> , \q<23> , \q<22> , \q<21> , 
        \q<20> , \q<19> , \q<18> , \q<17> , \q<16> , \q<15> , \q<14> , \q<13> , 
        \q<12> , \q<11> , \q<10> , \q<9> , \q<8> , \q<7> , \q<6> , \q<5> , 
        \q<4> , \q<3> , \q<2> , \q<1> , \q<0> }) );
  input clk, reset, \d<31> , \d<30> , \d<29> , \d<28> , \d<27> , \d<26> ,
         \d<25> , \d<24> , \d<23> , \d<22> , \d<21> , \d<20> , \d<19> ,
         \d<18> , \d<17> , \d<16> , \d<15> , \d<14> , \d<13> , \d<12> ,
         \d<11> , \d<10> , \d<9> , \d<8> , \d<7> , \d<6> , \d<5> , \d<4> ,
         \d<3> , \d<2> , \d<1> , \d<0> ;
  output \q<31> , \q<30> , \q<29> , \q<28> , \q<27> , \q<26> , \q<25> ,
         \q<24> , \q<23> , \q<22> , \q<21> , \q<20> , \q<19> , \q<18> ,
         \q<17> , \q<16> , \q<15> , \q<14> , \q<13> , \q<12> , \q<11> ,
         \q<10> , \q<9> , \q<8> , \q<7> , \q<6> , \q<5> , \q<4> , \q<3> ,
         \q<2> , \q<1> , \q<0> ;
  wire   n25, n26, n27, n28;

  DFFRHQX1 \q_reg<1>  ( .D(\d<1> ), .CK(clk), .RN(n25), .Q(\q<1> ) );
  DFFRHQX1 \q_reg<0>  ( .D(\d<0> ), .CK(clk), .RN(n26), .Q(\q<0> ) );
  DFFRHQX1 \q_reg<31>  ( .D(\d<31> ), .CK(clk), .RN(n25), .Q(\q<31> ) );
  DFFRHQX1 \q_reg<30>  ( .D(\d<30> ), .CK(clk), .RN(n26), .Q(\q<30> ) );
  DFFRHQX1 \q_reg<29>  ( .D(\d<29> ), .CK(clk), .RN(n25), .Q(\q<29> ) );
  DFFRHQX1 \q_reg<28>  ( .D(\d<28> ), .CK(clk), .RN(n26), .Q(\q<28> ) );
  DFFRHQX1 \q_reg<27>  ( .D(\d<27> ), .CK(clk), .RN(n28), .Q(\q<27> ) );
  DFFRHQX1 \q_reg<26>  ( .D(\d<26> ), .CK(clk), .RN(n28), .Q(\q<26> ) );
  DFFRHQX1 \q_reg<25>  ( .D(\d<25> ), .CK(clk), .RN(n26), .Q(\q<25> ) );
  DFFRHQX1 \q_reg<24>  ( .D(\d<24> ), .CK(clk), .RN(n26), .Q(\q<24> ) );
  DFFRHQX1 \q_reg<23>  ( .D(\d<23> ), .CK(clk), .RN(n26), .Q(\q<23> ) );
  DFFRHQX1 \q_reg<22>  ( .D(\d<22> ), .CK(clk), .RN(n26), .Q(\q<22> ) );
  DFFRHQX1 \q_reg<21>  ( .D(\d<21> ), .CK(clk), .RN(n26), .Q(\q<21> ) );
  DFFRHQX1 \q_reg<20>  ( .D(\d<20> ), .CK(clk), .RN(n26), .Q(\q<20> ) );
  DFFRHQX1 \q_reg<19>  ( .D(\d<19> ), .CK(clk), .RN(n26), .Q(\q<19> ) );
  DFFRHQX1 \q_reg<18>  ( .D(\d<18> ), .CK(clk), .RN(n26), .Q(\q<18> ) );
  DFFRHQX1 \q_reg<17>  ( .D(\d<17> ), .CK(clk), .RN(n26), .Q(\q<17> ) );
  DFFRHQX1 \q_reg<16>  ( .D(\d<16> ), .CK(clk), .RN(n26), .Q(\q<16> ) );
  DFFRHQX1 \q_reg<15>  ( .D(\d<15> ), .CK(clk), .RN(n26), .Q(\q<15> ) );
  DFFRHQX1 \q_reg<14>  ( .D(\d<14> ), .CK(clk), .RN(n26), .Q(\q<14> ) );
  DFFRHQX1 \q_reg<13>  ( .D(\d<13> ), .CK(clk), .RN(n25), .Q(\q<13> ) );
  DFFRHQX1 \q_reg<12>  ( .D(\d<12> ), .CK(clk), .RN(n25), .Q(\q<12> ) );
  DFFRHQX1 \q_reg<11>  ( .D(\d<11> ), .CK(clk), .RN(n25), .Q(\q<11> ) );
  DFFRHQX1 \q_reg<10>  ( .D(\d<10> ), .CK(clk), .RN(n25), .Q(\q<10> ) );
  DFFRHQX1 \q_reg<9>  ( .D(\d<9> ), .CK(clk), .RN(n25), .Q(\q<9> ) );
  DFFRHQX1 \q_reg<8>  ( .D(\d<8> ), .CK(clk), .RN(n25), .Q(\q<8> ) );
  DFFRHQX1 \q_reg<7>  ( .D(\d<7> ), .CK(clk), .RN(n25), .Q(\q<7> ) );
  DFFRHQX1 \q_reg<6>  ( .D(\d<6> ), .CK(clk), .RN(n25), .Q(\q<6> ) );
  DFFRHQX1 \q_reg<5>  ( .D(\d<5> ), .CK(clk), .RN(n25), .Q(\q<5> ) );
  DFFRHQX1 \q_reg<4>  ( .D(\d<4> ), .CK(clk), .RN(n25), .Q(\q<4> ) );
  DFFRHQX1 \q_reg<3>  ( .D(\d<3> ), .CK(clk), .RN(n25), .Q(\q<3> ) );
  DFFRHQX1 \q_reg<2>  ( .D(\d<2> ), .CK(clk), .RN(n25), .Q(\q<2> ) );
  CLKINVX3 U3 ( .A(n27), .Y(n26) );
  CLKINVX3 U4 ( .A(n27), .Y(n25) );
  INVX1 U5 ( .A(n28), .Y(n27) );
  INVXL U6 ( .A(reset), .Y(n28) );
endmodule


module flopr_WIDTH32_3 ( clk, reset, .d({\d<31> , \d<30> , \d<29> , \d<28> , 
        \d<27> , \d<26> , \d<25> , \d<24> , \d<23> , \d<22> , \d<21> , \d<20> , 
        \d<19> , \d<18> , \d<17> , \d<16> , \d<15> , \d<14> , \d<13> , \d<12> , 
        \d<11> , \d<10> , \d<9> , \d<8> , \d<7> , \d<6> , \d<5> , \d<4> , 
        \d<3> , \d<2> , \d<1> , \d<0> }), .q({\q<31> , \q<30> , \q<29> , 
        \q<28> , \q<27> , \q<26> , \q<25> , \q<24> , \q<23> , \q<22> , \q<21> , 
        \q<20> , \q<19> , \q<18> , \q<17> , \q<16> , \q<15> , \q<14> , \q<13> , 
        \q<12> , \q<11> , \q<10> , \q<9> , \q<8> , \q<7> , \q<6> , \q<5> , 
        \q<4> , \q<3> , \q<2> , \q<1> , \q<0> }) );
  input clk, reset, \d<31> , \d<30> , \d<29> , \d<28> , \d<27> , \d<26> ,
         \d<25> , \d<24> , \d<23> , \d<22> , \d<21> , \d<20> , \d<19> ,
         \d<18> , \d<17> , \d<16> , \d<15> , \d<14> , \d<13> , \d<12> ,
         \d<11> , \d<10> , \d<9> , \d<8> , \d<7> , \d<6> , \d<5> , \d<4> ,
         \d<3> , \d<2> , \d<1> , \d<0> ;
  output \q<31> , \q<30> , \q<29> , \q<28> , \q<27> , \q<26> , \q<25> ,
         \q<24> , \q<23> , \q<22> , \q<21> , \q<20> , \q<19> , \q<18> ,
         \q<17> , \q<16> , \q<15> , \q<14> , \q<13> , \q<12> , \q<11> ,
         \q<10> , \q<9> , \q<8> , \q<7> , \q<6> , \q<5> , \q<4> , \q<3> ,
         \q<2> , \q<1> , \q<0> ;
  wire   n25, n26, n27, n28;

  DFFRHQX1 \q_reg<31>  ( .D(\d<31> ), .CK(clk), .RN(n25), .Q(\q<31> ) );
  DFFRHQX1 \q_reg<30>  ( .D(\d<30> ), .CK(clk), .RN(n26), .Q(\q<30> ) );
  DFFRHQX1 \q_reg<29>  ( .D(\d<29> ), .CK(clk), .RN(n25), .Q(\q<29> ) );
  DFFRHQX1 \q_reg<28>  ( .D(\d<28> ), .CK(clk), .RN(n26), .Q(\q<28> ) );
  DFFRHQX1 \q_reg<27>  ( .D(\d<27> ), .CK(clk), .RN(n25), .Q(\q<27> ) );
  DFFRHQX1 \q_reg<26>  ( .D(\d<26> ), .CK(clk), .RN(n26), .Q(\q<26> ) );
  DFFRHQX1 \q_reg<25>  ( .D(\d<25> ), .CK(clk), .RN(n28), .Q(\q<25> ) );
  DFFRHQX1 \q_reg<24>  ( .D(\d<24> ), .CK(clk), .RN(n28), .Q(\q<24> ) );
  DFFRHQX1 \q_reg<23>  ( .D(\d<23> ), .CK(clk), .RN(n26), .Q(\q<23> ) );
  DFFRHQX1 \q_reg<22>  ( .D(\d<22> ), .CK(clk), .RN(n26), .Q(\q<22> ) );
  DFFRHQX1 \q_reg<21>  ( .D(\d<21> ), .CK(clk), .RN(n26), .Q(\q<21> ) );
  DFFRHQX1 \q_reg<20>  ( .D(\d<20> ), .CK(clk), .RN(n26), .Q(\q<20> ) );
  DFFRHQX1 \q_reg<19>  ( .D(\d<19> ), .CK(clk), .RN(n26), .Q(\q<19> ) );
  DFFRHQX1 \q_reg<18>  ( .D(\d<18> ), .CK(clk), .RN(n26), .Q(\q<18> ) );
  DFFRHQX1 \q_reg<17>  ( .D(\d<17> ), .CK(clk), .RN(n26), .Q(\q<17> ) );
  DFFRHQX1 \q_reg<16>  ( .D(\d<16> ), .CK(clk), .RN(n26), .Q(\q<16> ) );
  DFFRHQX1 \q_reg<15>  ( .D(\d<15> ), .CK(clk), .RN(n26), .Q(\q<15> ) );
  DFFRHQX1 \q_reg<14>  ( .D(\d<14> ), .CK(clk), .RN(n26), .Q(\q<14> ) );
  DFFRHQX1 \q_reg<13>  ( .D(\d<13> ), .CK(clk), .RN(n26), .Q(\q<13> ) );
  DFFRHQX1 \q_reg<12>  ( .D(\d<12> ), .CK(clk), .RN(n26), .Q(\q<12> ) );
  DFFRHQX1 \q_reg<11>  ( .D(\d<11> ), .CK(clk), .RN(n25), .Q(\q<11> ) );
  DFFRHQX1 \q_reg<10>  ( .D(\d<10> ), .CK(clk), .RN(n25), .Q(\q<10> ) );
  DFFRHQX1 \q_reg<9>  ( .D(\d<9> ), .CK(clk), .RN(n25), .Q(\q<9> ) );
  DFFRHQX1 \q_reg<8>  ( .D(\d<8> ), .CK(clk), .RN(n25), .Q(\q<8> ) );
  DFFRHQX1 \q_reg<7>  ( .D(\d<7> ), .CK(clk), .RN(n25), .Q(\q<7> ) );
  DFFRHQX1 \q_reg<6>  ( .D(\d<6> ), .CK(clk), .RN(n25), .Q(\q<6> ) );
  DFFRHQX1 \q_reg<5>  ( .D(\d<5> ), .CK(clk), .RN(n25), .Q(\q<5> ) );
  DFFRHQX1 \q_reg<4>  ( .D(\d<4> ), .CK(clk), .RN(n25), .Q(\q<4> ) );
  DFFRHQX1 \q_reg<3>  ( .D(\d<3> ), .CK(clk), .RN(n25), .Q(\q<3> ) );
  DFFRHQX1 \q_reg<2>  ( .D(\d<2> ), .CK(clk), .RN(n25), .Q(\q<2> ) );
  DFFRHQX1 \q_reg<1>  ( .D(\d<1> ), .CK(clk), .RN(n25), .Q(\q<1> ) );
  DFFRHQX1 \q_reg<0>  ( .D(\d<0> ), .CK(clk), .RN(n25), .Q(\q<0> ) );
  CLKINVX3 U3 ( .A(n27), .Y(n26) );
  CLKINVX3 U4 ( .A(n27), .Y(n25) );
  INVX1 U5 ( .A(n28), .Y(n27) );
  INVXL U6 ( .A(reset), .Y(n28) );
endmodule


module flopr_WIDTH32_2 ( clk, reset, .d({\d<31> , \d<30> , \d<29> , \d<28> , 
        \d<27> , \d<26> , \d<25> , \d<24> , \d<23> , \d<22> , \d<21> , \d<20> , 
        \d<19> , \d<18> , \d<17> , \d<16> , \d<15> , \d<14> , \d<13> , \d<12> , 
        \d<11> , \d<10> , \d<9> , \d<8> , \d<7> , \d<6> , \d<5> , \d<4> , 
        \d<3> , \d<2> , \d<1> , \d<0> }), .q({\q<31> , \q<30> , \q<29> , 
        \q<28> , \q<27> , \q<26> , \q<25> , \q<24> , \q<23> , \q<22> , \q<21> , 
        \q<20> , \q<19> , \q<18> , \q<17> , \q<16> , \q<15> , \q<14> , \q<13> , 
        \q<12> , \q<11> , \q<10> , \q<9> , \q<8> , \q<7> , \q<6> , \q<5> , 
        \q<4> , \q<3> , \q<2> , \q<1> , \q<0> }) );
  input clk, reset, \d<31> , \d<30> , \d<29> , \d<28> , \d<27> , \d<26> ,
         \d<25> , \d<24> , \d<23> , \d<22> , \d<21> , \d<20> , \d<19> ,
         \d<18> , \d<17> , \d<16> , \d<15> , \d<14> , \d<13> , \d<12> ,
         \d<11> , \d<10> , \d<9> , \d<8> , \d<7> , \d<6> , \d<5> , \d<4> ,
         \d<3> , \d<2> , \d<1> , \d<0> ;
  output \q<31> , \q<30> , \q<29> , \q<28> , \q<27> , \q<26> , \q<25> ,
         \q<24> , \q<23> , \q<22> , \q<21> , \q<20> , \q<19> , \q<18> ,
         \q<17> , \q<16> , \q<15> , \q<14> , \q<13> , \q<12> , \q<11> ,
         \q<10> , \q<9> , \q<8> , \q<7> , \q<6> , \q<5> , \q<4> , \q<3> ,
         \q<2> , \q<1> , \q<0> ;
  wire   n25, n26, n27, n28;

  DFFRHQX1 \q_reg<31>  ( .D(\d<31> ), .CK(clk), .RN(n25), .Q(\q<31> ) );
  DFFRHQX1 \q_reg<30>  ( .D(\d<30> ), .CK(clk), .RN(n26), .Q(\q<30> ) );
  DFFRHQX1 \q_reg<29>  ( .D(\d<29> ), .CK(clk), .RN(n25), .Q(\q<29> ) );
  DFFRHQX1 \q_reg<28>  ( .D(\d<28> ), .CK(clk), .RN(n26), .Q(\q<28> ) );
  DFFRHQX1 \q_reg<27>  ( .D(\d<27> ), .CK(clk), .RN(n25), .Q(\q<27> ) );
  DFFRHQX1 \q_reg<26>  ( .D(\d<26> ), .CK(clk), .RN(n26), .Q(\q<26> ) );
  DFFRHQX1 \q_reg<25>  ( .D(\d<25> ), .CK(clk), .RN(n28), .Q(\q<25> ) );
  DFFRHQX1 \q_reg<24>  ( .D(\d<24> ), .CK(clk), .RN(n28), .Q(\q<24> ) );
  DFFRHQX1 \q_reg<23>  ( .D(\d<23> ), .CK(clk), .RN(n26), .Q(\q<23> ) );
  DFFRHQX1 \q_reg<22>  ( .D(\d<22> ), .CK(clk), .RN(n26), .Q(\q<22> ) );
  DFFRHQX1 \q_reg<21>  ( .D(\d<21> ), .CK(clk), .RN(n26), .Q(\q<21> ) );
  DFFRHQX1 \q_reg<20>  ( .D(\d<20> ), .CK(clk), .RN(n26), .Q(\q<20> ) );
  DFFRHQX1 \q_reg<19>  ( .D(\d<19> ), .CK(clk), .RN(n26), .Q(\q<19> ) );
  DFFRHQX1 \q_reg<18>  ( .D(\d<18> ), .CK(clk), .RN(n26), .Q(\q<18> ) );
  DFFRHQX1 \q_reg<17>  ( .D(\d<17> ), .CK(clk), .RN(n26), .Q(\q<17> ) );
  DFFRHQX1 \q_reg<16>  ( .D(\d<16> ), .CK(clk), .RN(n26), .Q(\q<16> ) );
  DFFRHQX1 \q_reg<15>  ( .D(\d<15> ), .CK(clk), .RN(n26), .Q(\q<15> ) );
  DFFRHQX1 \q_reg<14>  ( .D(\d<14> ), .CK(clk), .RN(n26), .Q(\q<14> ) );
  DFFRHQX1 \q_reg<13>  ( .D(\d<13> ), .CK(clk), .RN(n26), .Q(\q<13> ) );
  DFFRHQX1 \q_reg<12>  ( .D(\d<12> ), .CK(clk), .RN(n26), .Q(\q<12> ) );
  DFFRHQX1 \q_reg<11>  ( .D(\d<11> ), .CK(clk), .RN(n25), .Q(\q<11> ) );
  DFFRHQX1 \q_reg<10>  ( .D(\d<10> ), .CK(clk), .RN(n25), .Q(\q<10> ) );
  DFFRHQX1 \q_reg<9>  ( .D(\d<9> ), .CK(clk), .RN(n25), .Q(\q<9> ) );
  DFFRHQX1 \q_reg<8>  ( .D(\d<8> ), .CK(clk), .RN(n25), .Q(\q<8> ) );
  DFFRHQX1 \q_reg<7>  ( .D(\d<7> ), .CK(clk), .RN(n25), .Q(\q<7> ) );
  DFFRHQX1 \q_reg<6>  ( .D(\d<6> ), .CK(clk), .RN(n25), .Q(\q<6> ) );
  DFFRHQX1 \q_reg<5>  ( .D(\d<5> ), .CK(clk), .RN(n25), .Q(\q<5> ) );
  DFFRHQX1 \q_reg<4>  ( .D(\d<4> ), .CK(clk), .RN(n25), .Q(\q<4> ) );
  DFFRHQX1 \q_reg<3>  ( .D(\d<3> ), .CK(clk), .RN(n25), .Q(\q<3> ) );
  DFFRHQX1 \q_reg<2>  ( .D(\d<2> ), .CK(clk), .RN(n25), .Q(\q<2> ) );
  DFFRHQX1 \q_reg<1>  ( .D(\d<1> ), .CK(clk), .RN(n25), .Q(\q<1> ) );
  DFFRHQX1 \q_reg<0>  ( .D(\d<0> ), .CK(clk), .RN(n25), .Q(\q<0> ) );
  CLKINVX3 U3 ( .A(n27), .Y(n26) );
  CLKINVX3 U4 ( .A(n27), .Y(n25) );
  INVX1 U5 ( .A(n28), .Y(n27) );
  INVXL U6 ( .A(reset), .Y(n28) );
endmodule


module flopr_WIDTH32_1 ( clk, reset, .d({\d<31> , \d<30> , \d<29> , \d<28> , 
        \d<27> , \d<26> , \d<25> , \d<24> , \d<23> , \d<22> , \d<21> , \d<20> , 
        \d<19> , \d<18> , \d<17> , \d<16> , \d<15> , \d<14> , \d<13> , \d<12> , 
        \d<11> , \d<10> , \d<9> , \d<8> , \d<7> , \d<6> , \d<5> , \d<4> , 
        \d<3> , \d<2> , \d<1> , \d<0> }), .q({\q<31> , \q<30> , \q<29> , 
        \q<28> , \q<27> , \q<26> , \q<25> , \q<24> , \q<23> , \q<22> , \q<21> , 
        \q<20> , \q<19> , \q<18> , \q<17> , \q<16> , \q<15> , \q<14> , \q<13> , 
        \q<12> , \q<11> , \q<10> , \q<9> , \q<8> , \q<7> , \q<6> , \q<5> , 
        \q<4> , \q<3> , \q<2> , \q<1> , \q<0> }) );
  input clk, reset, \d<31> , \d<30> , \d<29> , \d<28> , \d<27> , \d<26> ,
         \d<25> , \d<24> , \d<23> , \d<22> , \d<21> , \d<20> , \d<19> ,
         \d<18> , \d<17> , \d<16> , \d<15> , \d<14> , \d<13> , \d<12> ,
         \d<11> , \d<10> , \d<9> , \d<8> , \d<7> , \d<6> , \d<5> , \d<4> ,
         \d<3> , \d<2> , \d<1> , \d<0> ;
  output \q<31> , \q<30> , \q<29> , \q<28> , \q<27> , \q<26> , \q<25> ,
         \q<24> , \q<23> , \q<22> , \q<21> , \q<20> , \q<19> , \q<18> ,
         \q<17> , \q<16> , \q<15> , \q<14> , \q<13> , \q<12> , \q<11> ,
         \q<10> , \q<9> , \q<8> , \q<7> , \q<6> , \q<5> , \q<4> , \q<3> ,
         \q<2> , \q<1> , \q<0> ;
  wire   n25, n26, n27, n28;

  DFFRHQX1 \q_reg<31>  ( .D(\d<31> ), .CK(clk), .RN(n25), .Q(\q<31> ) );
  DFFRHQX1 \q_reg<30>  ( .D(\d<30> ), .CK(clk), .RN(n26), .Q(\q<30> ) );
  DFFRHQX1 \q_reg<29>  ( .D(\d<29> ), .CK(clk), .RN(n25), .Q(\q<29> ) );
  DFFRHQX1 \q_reg<28>  ( .D(\d<28> ), .CK(clk), .RN(n26), .Q(\q<28> ) );
  DFFRHQX1 \q_reg<27>  ( .D(\d<27> ), .CK(clk), .RN(n25), .Q(\q<27> ) );
  DFFRHQX1 \q_reg<26>  ( .D(\d<26> ), .CK(clk), .RN(n26), .Q(\q<26> ) );
  DFFRHQX1 \q_reg<25>  ( .D(\d<25> ), .CK(clk), .RN(n28), .Q(\q<25> ) );
  DFFRHQX1 \q_reg<24>  ( .D(\d<24> ), .CK(clk), .RN(n28), .Q(\q<24> ) );
  DFFRHQX1 \q_reg<23>  ( .D(\d<23> ), .CK(clk), .RN(n26), .Q(\q<23> ) );
  DFFRHQX1 \q_reg<22>  ( .D(\d<22> ), .CK(clk), .RN(n26), .Q(\q<22> ) );
  DFFRHQX1 \q_reg<21>  ( .D(\d<21> ), .CK(clk), .RN(n26), .Q(\q<21> ) );
  DFFRHQX1 \q_reg<20>  ( .D(\d<20> ), .CK(clk), .RN(n26), .Q(\q<20> ) );
  DFFRHQX1 \q_reg<19>  ( .D(\d<19> ), .CK(clk), .RN(n26), .Q(\q<19> ) );
  DFFRHQX1 \q_reg<18>  ( .D(\d<18> ), .CK(clk), .RN(n26), .Q(\q<18> ) );
  DFFRHQX1 \q_reg<17>  ( .D(\d<17> ), .CK(clk), .RN(n26), .Q(\q<17> ) );
  DFFRHQX1 \q_reg<16>  ( .D(\d<16> ), .CK(clk), .RN(n26), .Q(\q<16> ) );
  DFFRHQX1 \q_reg<15>  ( .D(\d<15> ), .CK(clk), .RN(n26), .Q(\q<15> ) );
  DFFRHQX1 \q_reg<14>  ( .D(\d<14> ), .CK(clk), .RN(n26), .Q(\q<14> ) );
  DFFRHQX1 \q_reg<13>  ( .D(\d<13> ), .CK(clk), .RN(n26), .Q(\q<13> ) );
  DFFRHQX1 \q_reg<12>  ( .D(\d<12> ), .CK(clk), .RN(n26), .Q(\q<12> ) );
  DFFRHQX1 \q_reg<9>  ( .D(\d<9> ), .CK(clk), .RN(n25), .Q(\q<9> ) );
  DFFRHQX1 \q_reg<11>  ( .D(\d<11> ), .CK(clk), .RN(n25), .Q(\q<11> ) );
  DFFRHQX1 \q_reg<10>  ( .D(\d<10> ), .CK(clk), .RN(n25), .Q(\q<10> ) );
  DFFRHQX1 \q_reg<8>  ( .D(\d<8> ), .CK(clk), .RN(n25), .Q(\q<8> ) );
  DFFRHQX1 \q_reg<7>  ( .D(\d<7> ), .CK(clk), .RN(n25), .Q(\q<7> ) );
  DFFRHQX1 \q_reg<6>  ( .D(\d<6> ), .CK(clk), .RN(n25), .Q(\q<6> ) );
  DFFRHQX1 \q_reg<5>  ( .D(\d<5> ), .CK(clk), .RN(n25), .Q(\q<5> ) );
  DFFRHQX1 \q_reg<4>  ( .D(\d<4> ), .CK(clk), .RN(n25), .Q(\q<4> ) );
  DFFRHQX1 \q_reg<3>  ( .D(\d<3> ), .CK(clk), .RN(n25), .Q(\q<3> ) );
  DFFRHQX1 \q_reg<2>  ( .D(\d<2> ), .CK(clk), .RN(n25), .Q(\q<2> ) );
  DFFRHQX1 \q_reg<1>  ( .D(\d<1> ), .CK(clk), .RN(n25), .Q(\q<1> ) );
  DFFRHQX1 \q_reg<0>  ( .D(\d<0> ), .CK(clk), .RN(n25), .Q(\q<0> ) );
  CLKINVX3 U3 ( .A(n27), .Y(n26) );
  CLKINVX3 U4 ( .A(n27), .Y(n25) );
  INVX1 U5 ( .A(n28), .Y(n27) );
  INVXL U6 ( .A(reset), .Y(n28) );
endmodule


module mux2_WIDTH32 ( .d0({\d0<31> , \d0<30> , \d0<29> , \d0<28> , \d0<27> , 
        \d0<26> , \d0<25> , \d0<24> , \d0<23> , \d0<22> , \d0<21> , \d0<20> , 
        \d0<19> , \d0<18> , \d0<17> , \d0<16> , \d0<15> , \d0<14> , \d0<13> , 
        \d0<12> , \d0<11> , \d0<10> , \d0<9> , \d0<8> , \d0<7> , \d0<6> , 
        \d0<5> , \d0<4> , \d0<3> , \d0<2> , \d0<1> , \d0<0> }), .d1({\d1<31> , 
        \d1<30> , \d1<29> , \d1<28> , \d1<27> , \d1<26> , \d1<25> , \d1<24> , 
        \d1<23> , \d1<22> , \d1<21> , \d1<20> , \d1<19> , \d1<18> , \d1<17> , 
        \d1<16> , \d1<15> , \d1<14> , \d1<13> , \d1<12> , \d1<11> , \d1<10> , 
        \d1<9> , \d1<8> , \d1<7> , \d1<6> , \d1<5> , \d1<4> , \d1<3> , \d1<2> , 
        \d1<1> , \d1<0> }), s, .y({\y<31> , \y<30> , \y<29> , \y<28> , \y<27> , 
        \y<26> , \y<25> , \y<24> , \y<23> , \y<22> , \y<21> , \y<20> , \y<19> , 
        \y<18> , \y<17> , \y<16> , \y<15> , \y<14> , \y<13> , \y<12> , \y<11> , 
        \y<10> , \y<9> , \y<8> , \y<7> , \y<6> , \y<5> , \y<4> , \y<3> , 
        \y<2> , \y<1> , \y<0> }) );
  input \d0<31> , \d0<30> , \d0<29> , \d0<28> , \d0<27> , \d0<26> , \d0<25> ,
         \d0<24> , \d0<23> , \d0<22> , \d0<21> , \d0<20> , \d0<19> , \d0<18> ,
         \d0<17> , \d0<16> , \d0<15> , \d0<14> , \d0<13> , \d0<12> , \d0<11> ,
         \d0<10> , \d0<9> , \d0<8> , \d0<7> , \d0<6> , \d0<5> , \d0<4> ,
         \d0<3> , \d0<2> , \d0<1> , \d0<0> , \d1<31> , \d1<30> , \d1<29> ,
         \d1<28> , \d1<27> , \d1<26> , \d1<25> , \d1<24> , \d1<23> , \d1<22> ,
         \d1<21> , \d1<20> , \d1<19> , \d1<18> , \d1<17> , \d1<16> , \d1<15> ,
         \d1<14> , \d1<13> , \d1<12> , \d1<11> , \d1<10> , \d1<9> , \d1<8> ,
         \d1<7> , \d1<6> , \d1<5> , \d1<4> , \d1<3> , \d1<2> , \d1<1> ,
         \d1<0> , s;
  output \y<31> , \y<30> , \y<29> , \y<28> , \y<27> , \y<26> , \y<25> ,
         \y<24> , \y<23> , \y<22> , \y<21> , \y<20> , \y<19> , \y<18> ,
         \y<17> , \y<16> , \y<15> , \y<14> , \y<13> , \y<12> , \y<11> ,
         \y<10> , \y<9> , \y<8> , \y<7> , \y<6> , \y<5> , \y<4> , \y<3> ,
         \y<2> , \y<1> , \y<0> ;
  wire   n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61,
         n62, n63, n64, n65, n83, n84, n85, n86, n87, n88, n89, n90;

  CLKINVX3 U1 ( .A(n90), .Y(n84) );
  CLKINVX3 U2 ( .A(n90), .Y(n85) );
  INVX1 U3 ( .A(n83), .Y(n87) );
  INVX1 U4 ( .A(n84), .Y(n86) );
  INVX1 U5 ( .A(n84), .Y(n89) );
  INVX1 U6 ( .A(n83), .Y(n88) );
  INVX1 U7 ( .A(n83), .Y(n90) );
  INVX1 U8 ( .A(s), .Y(n83) );
  INVX1 U9 ( .A(n41), .Y(\y<31> ) );
  AOI22X1 U10 ( .A0(\d0<31> ), .A1(n84), .B0(\d1<31> ), .B1(n88), .Y(n41) );
  INVX1 U11 ( .A(n44), .Y(\y<29> ) );
  AOI22X1 U12 ( .A0(\d0<29> ), .A1(n85), .B0(\d1<29> ), .B1(n86), .Y(n44) );
  INVX1 U13 ( .A(n45), .Y(\y<28> ) );
  AOI22X1 U14 ( .A0(\d0<28> ), .A1(n85), .B0(\d1<28> ), .B1(s), .Y(n45) );
  INVX1 U15 ( .A(n42), .Y(\y<30> ) );
  AOI22X1 U16 ( .A0(\d0<30> ), .A1(n85), .B0(\d1<30> ), .B1(n89), .Y(n42) );
  INVX1 U17 ( .A(n46), .Y(\y<27> ) );
  AOI22X1 U18 ( .A0(\d0<27> ), .A1(n85), .B0(\d1<27> ), .B1(n86), .Y(n46) );
  INVX1 U19 ( .A(n47), .Y(\y<26> ) );
  AOI22X1 U20 ( .A0(\d0<26> ), .A1(n85), .B0(\d1<26> ), .B1(n86), .Y(n47) );
  INVX1 U21 ( .A(n50), .Y(\y<23> ) );
  AOI22X1 U22 ( .A0(\d0<23> ), .A1(n85), .B0(\d1<23> ), .B1(s), .Y(n50) );
  INVX1 U23 ( .A(n51), .Y(\y<22> ) );
  AOI22X1 U24 ( .A0(\d0<22> ), .A1(n85), .B0(\d1<22> ), .B1(n88), .Y(n51) );
  INVX1 U25 ( .A(n49), .Y(\y<24> ) );
  AOI22X1 U26 ( .A0(\d0<24> ), .A1(n85), .B0(\d1<24> ), .B1(n86), .Y(n49) );
  INVX1 U27 ( .A(n48), .Y(\y<25> ) );
  AOI22X1 U28 ( .A0(\d0<25> ), .A1(n85), .B0(\d1<25> ), .B1(n86), .Y(n48) );
  INVX1 U29 ( .A(n52), .Y(\y<21> ) );
  AOI22X1 U30 ( .A0(\d0<21> ), .A1(n85), .B0(\d1<21> ), .B1(n89), .Y(n52) );
  INVX1 U31 ( .A(n57), .Y(\y<17> ) );
  AOI22X1 U32 ( .A0(\d0<17> ), .A1(n84), .B0(\d1<17> ), .B1(n87), .Y(n57) );
  INVX1 U33 ( .A(n56), .Y(\y<18> ) );
  AOI22X1 U34 ( .A0(\d0<18> ), .A1(n84), .B0(\d1<18> ), .B1(n89), .Y(n56) );
  INVX1 U35 ( .A(n55), .Y(\y<19> ) );
  AOI22X1 U36 ( .A0(\d0<19> ), .A1(n84), .B0(\d1<19> ), .B1(n88), .Y(n55) );
  INVX1 U37 ( .A(n53), .Y(\y<20> ) );
  AOI22X1 U38 ( .A0(\d0<20> ), .A1(n85), .B0(\d1<20> ), .B1(s), .Y(n53) );
  INVX1 U39 ( .A(n58), .Y(\y<16> ) );
  AOI22X1 U40 ( .A0(\d0<16> ), .A1(n84), .B0(\d1<16> ), .B1(s), .Y(n58) );
  INVX1 U41 ( .A(n62), .Y(\y<12> ) );
  AOI22X1 U42 ( .A0(\d0<12> ), .A1(n84), .B0(\d1<12> ), .B1(n90), .Y(n62) );
  INVX1 U43 ( .A(n61), .Y(\y<13> ) );
  AOI22X1 U44 ( .A0(\d0<13> ), .A1(n84), .B0(\d1<13> ), .B1(n89), .Y(n61) );
  INVX1 U45 ( .A(n59), .Y(\y<15> ) );
  AOI22X1 U46 ( .A0(\d0<15> ), .A1(n84), .B0(\d1<15> ), .B1(n89), .Y(n59) );
  INVX1 U47 ( .A(n60), .Y(\y<14> ) );
  AOI22X1 U48 ( .A0(\d0<14> ), .A1(n84), .B0(\d1<14> ), .B1(n89), .Y(n60) );
  INVX1 U49 ( .A(n36), .Y(\y<7> ) );
  AOI22X1 U50 ( .A0(\d0<7> ), .A1(n84), .B0(\d1<7> ), .B1(n86), .Y(n36) );
  INVX1 U51 ( .A(n63), .Y(\y<11> ) );
  AOI22X1 U52 ( .A0(\d0<11> ), .A1(n84), .B0(\d1<11> ), .B1(n88), .Y(n63) );
  INVX1 U53 ( .A(n64), .Y(\y<10> ) );
  AOI22X1 U54 ( .A0(\d0<10> ), .A1(n84), .B0(\d1<10> ), .B1(n89), .Y(n64) );
  INVX1 U55 ( .A(n35), .Y(\y<8> ) );
  AOI22X1 U56 ( .A0(\d0<8> ), .A1(n84), .B0(\d1<8> ), .B1(n86), .Y(n35) );
  INVX1 U57 ( .A(n34), .Y(\y<9> ) );
  AOI22X1 U58 ( .A0(\d0<9> ), .A1(n84), .B0(n88), .B1(\d1<9> ), .Y(n34) );
  INVX1 U59 ( .A(n39), .Y(\y<4> ) );
  AOI22X1 U60 ( .A0(\d0<4> ), .A1(n83), .B0(\d1<4> ), .B1(n87), .Y(n39) );
  INVX1 U61 ( .A(n38), .Y(\y<5> ) );
  AOI22X1 U62 ( .A0(\d0<5> ), .A1(n83), .B0(\d1<5> ), .B1(n87), .Y(n38) );
  INVX1 U63 ( .A(n43), .Y(\y<2> ) );
  AOI22X1 U64 ( .A0(\d0<2> ), .A1(n85), .B0(\d1<2> ), .B1(n88), .Y(n43) );
  INVX1 U65 ( .A(n40), .Y(\y<3> ) );
  AOI22X1 U66 ( .A0(\d0<3> ), .A1(n83), .B0(\d1<3> ), .B1(n87), .Y(n40) );
  INVX1 U67 ( .A(n37), .Y(\y<6> ) );
  AOI22X1 U68 ( .A0(\d0<6> ), .A1(n84), .B0(\d1<6> ), .B1(n90), .Y(n37) );
  INVX1 U69 ( .A(n65), .Y(\y<0> ) );
  AOI22X1 U70 ( .A0(\d0<0> ), .A1(n84), .B0(\d1<0> ), .B1(n88), .Y(n65) );
  INVX1 U71 ( .A(n54), .Y(\y<1> ) );
  AOI22X1 U72 ( .A0(\d0<1> ), .A1(n84), .B0(\d1<1> ), .B1(s), .Y(n54) );
endmodule


module mux2_WIDTH4_0 ( .d0({\d0<3> , \d0<2> , \d0<1> , \d0<0> }), .d1({\d1<3> , 
        \d1<2> , \d1<1> , \d1<0> }), s, .y({\y<3> , \y<2> , \y<1> , \y<0> })
 );
  input \d0<3> , \d0<2> , \d0<1> , \d0<0> , \d1<3> , \d1<2> , \d1<1> , \d1<0> ,
         s;
  output \y<3> , \y<2> , \y<1> , \y<0> ;
  wire   n6, n7, n8, n9, n15;

  INVX1 U1 ( .A(s), .Y(n15) );
  INVX1 U2 ( .A(n8), .Y(\y<1> ) );
  AOI22X1 U3 ( .A0(\d0<1> ), .A1(n15), .B0(\d1<1> ), .B1(s), .Y(n8) );
  INVX1 U4 ( .A(n6), .Y(\y<3> ) );
  AOI22X1 U5 ( .A0(\d0<3> ), .A1(n15), .B0(s), .B1(\d1<3> ), .Y(n6) );
  INVX1 U6 ( .A(n7), .Y(\y<2> ) );
  AOI22X1 U7 ( .A0(\d0<2> ), .A1(n15), .B0(\d1<2> ), .B1(s), .Y(n7) );
  INVX1 U8 ( .A(n9), .Y(\y<0> ) );
  AOI22X1 U9 ( .A0(\d0<0> ), .A1(n15), .B0(\d1<0> ), .B1(s), .Y(n9) );
endmodule


module mux2_WIDTH4_1 ( .d0({\d0<3> , \d0<2> , \d0<1> , \d0<0> }), .d1({\d1<3> , 
        \d1<2> , \d1<1> , \d1<0> }), s, .y({\y<3> , \y<2> , \y<1> , \y<0> })
 );
  input \d0<3> , \d0<2> , \d0<1> , \d0<0> , \d1<3> , \d1<2> , \d1<1> , \d1<0> ,
         s;
  output \y<3> , \y<2> , \y<1> , \y<0> ;
  wire   n6, n7, n8, n9, n19;

  INVX1 U1 ( .A(n6), .Y(\y<3> ) );
  INVX1 U2 ( .A(s), .Y(n19) );
  AOI22X1 U3 ( .A0(\d0<3> ), .A1(n19), .B0(s), .B1(\d1<3> ), .Y(n6) );
  INVX1 U4 ( .A(n8), .Y(\y<1> ) );
  AOI22X1 U5 ( .A0(\d0<1> ), .A1(n19), .B0(\d1<1> ), .B1(s), .Y(n8) );
  INVX1 U6 ( .A(n7), .Y(\y<2> ) );
  AOI22X1 U7 ( .A0(\d0<2> ), .A1(n19), .B0(\d1<2> ), .B1(s), .Y(n7) );
  INVX1 U8 ( .A(n9), .Y(\y<0> ) );
  AOI22X1 U9 ( .A0(\d0<0> ), .A1(n19), .B0(\d1<0> ), .B1(s), .Y(n9) );
endmodule


module mux3_WIDTH32_0 ( .d0({\d0<31> , \d0<30> , \d0<29> , \d0<28> , \d0<27> , 
        \d0<26> , \d0<25> , \d0<24> , \d0<23> , \d0<22> , \d0<21> , \d0<20> , 
        \d0<19> , \d0<18> , \d0<17> , \d0<16> , \d0<15> , \d0<14> , \d0<13> , 
        \d0<12> , \d0<11> , \d0<10> , \d0<9> , \d0<8> , \d0<7> , \d0<6> , 
        \d0<5> , \d0<4> , \d0<3> , \d0<2> , \d0<1> , \d0<0> }), .d1({\d1<31> , 
        \d1<30> , \d1<29> , \d1<28> , \d1<27> , \d1<26> , \d1<25> , \d1<24> , 
        \d1<23> , \d1<22> , \d1<21> , \d1<20> , \d1<19> , \d1<18> , \d1<17> , 
        \d1<16> , \d1<15> , \d1<14> , \d1<13> , \d1<12> , \d1<11> , \d1<10> , 
        \d1<9> , \d1<8> , \d1<7> , \d1<6> , \d1<5> , \d1<4> , \d1<3> , \d1<2> , 
        \d1<1> , \d1<0> }), .d2({\d2<31> , \d2<30> , \d2<29> , \d2<28> , 
        \d2<27> , \d2<26> , \d2<25> , \d2<24> , \d2<23> , \d2<22> , \d2<21> , 
        \d2<20> , \d2<19> , \d2<18> , \d2<17> , \d2<16> , \d2<15> , \d2<14> , 
        \d2<13> , \d2<12> , \d2<11> , \d2<10> , \d2<9> , \d2<8> , \d2<7> , 
        \d2<6> , \d2<5> , \d2<4> , \d2<3> , \d2<2> , \d2<1> , \d2<0> }), .s({
        \s<1> , \s<0> }), .y({\y<31> , \y<30> , \y<29> , \y<28> , \y<27> , 
        \y<26> , \y<25> , \y<24> , \y<23> , \y<22> , \y<21> , \y<20> , \y<19> , 
        \y<18> , \y<17> , \y<16> , \y<15> , \y<14> , \y<13> , \y<12> , \y<11> , 
        \y<10> , \y<9> , \y<8> , \y<7> , \y<6> , \y<5> , \y<4> , \y<3> , 
        \y<2> , \y<1> , \y<0> }) );
  input \d0<31> , \d0<30> , \d0<29> , \d0<28> , \d0<27> , \d0<26> , \d0<25> ,
         \d0<24> , \d0<23> , \d0<22> , \d0<21> , \d0<20> , \d0<19> , \d0<18> ,
         \d0<17> , \d0<16> , \d0<15> , \d0<14> , \d0<13> , \d0<12> , \d0<11> ,
         \d0<10> , \d0<9> , \d0<8> , \d0<7> , \d0<6> , \d0<5> , \d0<4> ,
         \d0<3> , \d0<2> , \d0<1> , \d0<0> , \d1<31> , \d1<30> , \d1<29> ,
         \d1<28> , \d1<27> , \d1<26> , \d1<25> , \d1<24> , \d1<23> , \d1<22> ,
         \d1<21> , \d1<20> , \d1<19> , \d1<18> , \d1<17> , \d1<16> , \d1<15> ,
         \d1<14> , \d1<13> , \d1<12> , \d1<11> , \d1<10> , \d1<9> , \d1<8> ,
         \d1<7> , \d1<6> , \d1<5> , \d1<4> , \d1<3> , \d1<2> , \d1<1> ,
         \d1<0> , \d2<31> , \d2<30> , \d2<29> , \d2<28> , \d2<27> , \d2<26> ,
         \d2<25> , \d2<24> , \d2<23> , \d2<22> , \d2<21> , \d2<20> , \d2<19> ,
         \d2<18> , \d2<17> , \d2<16> , \d2<15> , \d2<14> , \d2<13> , \d2<12> ,
         \d2<11> , \d2<10> , \d2<9> , \d2<8> , \d2<7> , \d2<6> , \d2<5> ,
         \d2<4> , \d2<3> , \d2<2> , \d2<1> , \d2<0> , \s<1> , \s<0> ;
  output \y<31> , \y<30> , \y<29> , \y<28> , \y<27> , \y<26> , \y<25> ,
         \y<24> , \y<23> , \y<22> , \y<21> , \y<20> , \y<19> , \y<18> ,
         \y<17> , \y<16> , \y<15> , \y<14> , \y<13> , \y<12> , \y<11> ,
         \y<10> , \y<9> , \y<8> , \y<7> , \y<6> , \y<5> , \y<4> , \y<3> ,
         \y<2> , \y<1> , \y<0> ;
  wire   n1, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n88, n89, n90, n91, n92, n93, n94, n95, n96;

  OR2X2 U1 ( .A(n96), .B(\s<0> ), .Y(n88) );
  OAI2BB1X1 U2 ( .A0N(\d2<0> ), .A1N(n96), .B0(n34), .Y(\y<0> ) );
  OAI2BB1X1 U3 ( .A0N(\d2<31> ), .A1N(n96), .B0(n10), .Y(\y<31> ) );
  CLKINVX3 U4 ( .A(n88), .Y(n93) );
  CLKINVX3 U5 ( .A(n91), .Y(n90) );
  CLKINVX3 U6 ( .A(n91), .Y(n89) );
  INVX1 U7 ( .A(n3), .Y(n91) );
  CLKINVX3 U8 ( .A(n88), .Y(n92) );
  NOR2BX1 U9 ( .AN(\s<0> ), .B(n96), .Y(n3) );
  CLKINVX3 U10 ( .A(n95), .Y(n96) );
  INVX1 U11 ( .A(n95), .Y(n94) );
  INVX1 U12 ( .A(\s<1> ), .Y(n95) );
  OAI2BB1X1 U13 ( .A0N(\d2<1> ), .A1N(n96), .B0(n23), .Y(\y<1> ) );
  AOI22X1 U14 ( .A0(\d0<1> ), .A1(n92), .B0(\d1<1> ), .B1(n89), .Y(n23) );
  OAI2BB1X1 U15 ( .A0N(\d2<2> ), .A1N(n96), .B0(n12), .Y(\y<2> ) );
  AOI22X1 U16 ( .A0(\d0<2> ), .A1(n93), .B0(\d1<2> ), .B1(n90), .Y(n12) );
  OAI2BB1X1 U17 ( .A0N(\d2<3> ), .A1N(n96), .B0(n9), .Y(\y<3> ) );
  AOI22X1 U18 ( .A0(\d0<3> ), .A1(n93), .B0(\d1<3> ), .B1(n90), .Y(n9) );
  AOI22X1 U19 ( .A0(\d0<0> ), .A1(n92), .B0(\d1<0> ), .B1(n89), .Y(n34) );
  OAI2BB1X1 U20 ( .A0N(n96), .A1N(\d2<9> ), .B0(n1), .Y(\y<9> ) );
  AOI22X1 U21 ( .A0(\d0<9> ), .A1(n93), .B0(\d1<9> ), .B1(n90), .Y(n1) );
  OAI2BB1X1 U22 ( .A0N(\d2<5> ), .A1N(n96), .B0(n7), .Y(\y<5> ) );
  AOI22X1 U23 ( .A0(\d0<5> ), .A1(n93), .B0(\d1<5> ), .B1(n90), .Y(n7) );
  OAI2BB1X1 U24 ( .A0N(\d2<7> ), .A1N(n96), .B0(n5), .Y(\y<7> ) );
  AOI22X1 U25 ( .A0(\d0<7> ), .A1(n93), .B0(\d1<7> ), .B1(n90), .Y(n5) );
  OAI2BB1X1 U26 ( .A0N(\d2<4> ), .A1N(n96), .B0(n8), .Y(\y<4> ) );
  AOI22X1 U27 ( .A0(\d0<4> ), .A1(n93), .B0(\d1<4> ), .B1(n90), .Y(n8) );
  OAI2BB1X1 U28 ( .A0N(\d2<6> ), .A1N(n96), .B0(n6), .Y(\y<6> ) );
  AOI22X1 U29 ( .A0(\d0<6> ), .A1(n93), .B0(\d1<6> ), .B1(n90), .Y(n6) );
  OAI2BB1X1 U30 ( .A0N(\d2<8> ), .A1N(n96), .B0(n4), .Y(\y<8> ) );
  AOI22X1 U31 ( .A0(\d0<8> ), .A1(n93), .B0(\d1<8> ), .B1(n90), .Y(n4) );
  OAI2BB1X1 U32 ( .A0N(\d2<10> ), .A1N(n96), .B0(n33), .Y(\y<10> ) );
  AOI22X1 U33 ( .A0(\d0<10> ), .A1(n92), .B0(\d1<10> ), .B1(n89), .Y(n33) );
  OAI2BB1X1 U34 ( .A0N(\d2<11> ), .A1N(n94), .B0(n32), .Y(\y<11> ) );
  AOI22X1 U35 ( .A0(\d0<11> ), .A1(n92), .B0(\d1<11> ), .B1(n89), .Y(n32) );
  OAI2BB1X1 U36 ( .A0N(\d2<12> ), .A1N(\s<1> ), .B0(n31), .Y(\y<12> ) );
  AOI22X1 U37 ( .A0(\d0<12> ), .A1(n92), .B0(\d1<12> ), .B1(n89), .Y(n31) );
  OAI2BB1X1 U38 ( .A0N(\d2<13> ), .A1N(\s<1> ), .B0(n30), .Y(\y<13> ) );
  AOI22X1 U39 ( .A0(\d0<13> ), .A1(n92), .B0(\d1<13> ), .B1(n89), .Y(n30) );
  OAI2BB1X1 U40 ( .A0N(\d2<14> ), .A1N(\s<1> ), .B0(n29), .Y(\y<14> ) );
  AOI22X1 U41 ( .A0(\d0<14> ), .A1(n92), .B0(\d1<14> ), .B1(n89), .Y(n29) );
  OAI2BB1X1 U42 ( .A0N(\d2<15> ), .A1N(\s<1> ), .B0(n28), .Y(\y<15> ) );
  AOI22X1 U43 ( .A0(\d0<15> ), .A1(n92), .B0(\d1<15> ), .B1(n89), .Y(n28) );
  OAI2BB1X1 U44 ( .A0N(\d2<16> ), .A1N(\s<1> ), .B0(n27), .Y(\y<16> ) );
  AOI22X1 U45 ( .A0(\d0<16> ), .A1(n92), .B0(\d1<16> ), .B1(n89), .Y(n27) );
  OAI2BB1X1 U46 ( .A0N(\d2<17> ), .A1N(\s<1> ), .B0(n26), .Y(\y<17> ) );
  AOI22X1 U47 ( .A0(\d0<17> ), .A1(n92), .B0(\d1<17> ), .B1(n89), .Y(n26) );
  OAI2BB1X1 U48 ( .A0N(\d2<18> ), .A1N(n94), .B0(n25), .Y(\y<18> ) );
  AOI22X1 U49 ( .A0(\d0<18> ), .A1(n92), .B0(\d1<18> ), .B1(n89), .Y(n25) );
  OAI2BB1X1 U50 ( .A0N(\d2<19> ), .A1N(n94), .B0(n24), .Y(\y<19> ) );
  AOI22X1 U51 ( .A0(\d0<19> ), .A1(n92), .B0(\d1<19> ), .B1(n89), .Y(n24) );
  OAI2BB1X1 U52 ( .A0N(\d2<20> ), .A1N(n94), .B0(n22), .Y(\y<20> ) );
  AOI22X1 U53 ( .A0(\d0<20> ), .A1(n93), .B0(\d1<20> ), .B1(n90), .Y(n22) );
  OAI2BB1X1 U54 ( .A0N(\d2<21> ), .A1N(n94), .B0(n21), .Y(\y<21> ) );
  AOI22X1 U55 ( .A0(\d0<21> ), .A1(n93), .B0(\d1<21> ), .B1(n90), .Y(n21) );
  OAI2BB1X1 U56 ( .A0N(\d2<22> ), .A1N(n94), .B0(n20), .Y(\y<22> ) );
  AOI22X1 U57 ( .A0(\d0<22> ), .A1(n93), .B0(\d1<22> ), .B1(n90), .Y(n20) );
  OAI2BB1X1 U58 ( .A0N(\d2<23> ), .A1N(n96), .B0(n19), .Y(\y<23> ) );
  AOI22X1 U59 ( .A0(\d0<23> ), .A1(n93), .B0(\d1<23> ), .B1(n90), .Y(n19) );
  OAI2BB1X1 U60 ( .A0N(\d2<24> ), .A1N(n96), .B0(n18), .Y(\y<24> ) );
  AOI22X1 U61 ( .A0(\d0<24> ), .A1(n93), .B0(\d1<24> ), .B1(n90), .Y(n18) );
  OAI2BB1X1 U62 ( .A0N(\d2<25> ), .A1N(n96), .B0(n17), .Y(\y<25> ) );
  AOI22X1 U63 ( .A0(\d0<25> ), .A1(n93), .B0(\d1<25> ), .B1(n90), .Y(n17) );
  OAI2BB1X1 U64 ( .A0N(\d2<26> ), .A1N(n96), .B0(n16), .Y(\y<26> ) );
  AOI22X1 U65 ( .A0(\d0<26> ), .A1(n93), .B0(\d1<26> ), .B1(n90), .Y(n16) );
  OAI2BB1X1 U66 ( .A0N(\d2<27> ), .A1N(n96), .B0(n15), .Y(\y<27> ) );
  AOI22X1 U67 ( .A0(\d0<27> ), .A1(n93), .B0(\d1<27> ), .B1(n90), .Y(n15) );
  OAI2BB1X1 U68 ( .A0N(\d2<28> ), .A1N(n96), .B0(n14), .Y(\y<28> ) );
  AOI22X1 U69 ( .A0(\d0<28> ), .A1(n93), .B0(\d1<28> ), .B1(n90), .Y(n14) );
  OAI2BB1X1 U70 ( .A0N(\d2<29> ), .A1N(n96), .B0(n13), .Y(\y<29> ) );
  AOI22X1 U71 ( .A0(\d0<29> ), .A1(n93), .B0(\d1<29> ), .B1(n90), .Y(n13) );
  AOI22X1 U72 ( .A0(\d0<31> ), .A1(n93), .B0(\d1<31> ), .B1(n90), .Y(n10) );
  OAI2BB1X1 U73 ( .A0N(\d2<30> ), .A1N(n96), .B0(n11), .Y(\y<30> ) );
  AOI22X1 U74 ( .A0(\d0<30> ), .A1(n93), .B0(\d1<30> ), .B1(n90), .Y(n11) );
endmodule


module mux3_WIDTH32_2 ( .d0({\d0<31> , \d0<30> , \d0<29> , \d0<28> , \d0<27> , 
        \d0<26> , \d0<25> , \d0<24> , \d0<23> , \d0<22> , \d0<21> , \d0<20> , 
        \d0<19> , \d0<18> , \d0<17> , \d0<16> , \d0<15> , \d0<14> , \d0<13> , 
        \d0<12> , \d0<11> , \d0<10> , \d0<9> , \d0<8> , \d0<7> , \d0<6> , 
        \d0<5> , \d0<4> , \d0<3> , \d0<2> , \d0<1> , \d0<0> }), .d1({\d1<31> , 
        \d1<30> , \d1<29> , \d1<28> , \d1<27> , \d1<26> , \d1<25> , \d1<24> , 
        \d1<23> , \d1<22> , \d1<21> , \d1<20> , \d1<19> , \d1<18> , \d1<17> , 
        \d1<16> , \d1<15> , \d1<14> , \d1<13> , \d1<12> , \d1<11> , \d1<10> , 
        \d1<9> , \d1<8> , \d1<7> , \d1<6> , \d1<5> , \d1<4> , \d1<3> , \d1<2> , 
        \d1<1> , \d1<0> }), .d2({\d2<31> , \d2<30> , \d2<29> , \d2<28> , 
        \d2<27> , \d2<26> , \d2<25> , \d2<24> , \d2<23> , \d2<22> , \d2<21> , 
        \d2<20> , \d2<19> , \d2<18> , \d2<17> , \d2<16> , \d2<15> , \d2<14> , 
        \d2<13> , \d2<12> , \d2<11> , \d2<10> , \d2<9> , \d2<8> , \d2<7> , 
        \d2<6> , \d2<5> , \d2<4> , \d2<3> , \d2<2> , \d2<1> , \d2<0> }), .s({
        \s<1> , \s<0> }), .y({\y<31> , \y<30> , \y<29> , \y<28> , \y<27> , 
        \y<26> , \y<25> , \y<24> , \y<23> , \y<22> , \y<21> , \y<20> , \y<19> , 
        \y<18> , \y<17> , \y<16> , \y<15> , \y<14> , \y<13> , \y<12> , \y<11> , 
        \y<10> , \y<9> , \y<8> , \y<7> , \y<6> , \y<5> , \y<4> , \y<3> , 
        \y<2> , \y<1> , \y<0> }) );
  input \d0<31> , \d0<30> , \d0<29> , \d0<28> , \d0<27> , \d0<26> , \d0<25> ,
         \d0<24> , \d0<23> , \d0<22> , \d0<21> , \d0<20> , \d0<19> , \d0<18> ,
         \d0<17> , \d0<16> , \d0<15> , \d0<14> , \d0<13> , \d0<12> , \d0<11> ,
         \d0<10> , \d0<9> , \d0<8> , \d0<7> , \d0<6> , \d0<5> , \d0<4> ,
         \d0<3> , \d0<2> , \d0<1> , \d0<0> , \d1<31> , \d1<30> , \d1<29> ,
         \d1<28> , \d1<27> , \d1<26> , \d1<25> , \d1<24> , \d1<23> , \d1<22> ,
         \d1<21> , \d1<20> , \d1<19> , \d1<18> , \d1<17> , \d1<16> , \d1<15> ,
         \d1<14> , \d1<13> , \d1<12> , \d1<11> , \d1<10> , \d1<9> , \d1<8> ,
         \d1<7> , \d1<6> , \d1<5> , \d1<4> , \d1<3> , \d1<2> , \d1<1> ,
         \d1<0> , \d2<31> , \d2<30> , \d2<29> , \d2<28> , \d2<27> , \d2<26> ,
         \d2<25> , \d2<24> , \d2<23> , \d2<22> , \d2<21> , \d2<20> , \d2<19> ,
         \d2<18> , \d2<17> , \d2<16> , \d2<15> , \d2<14> , \d2<13> , \d2<12> ,
         \d2<11> , \d2<10> , \d2<9> , \d2<8> , \d2<7> , \d2<6> , \d2<5> ,
         \d2<4> , \d2<3> , \d2<2> , \d2<1> , \d2<0> , \s<1> , \s<0> ;
  output \y<31> , \y<30> , \y<29> , \y<28> , \y<27> , \y<26> , \y<25> ,
         \y<24> , \y<23> , \y<22> , \y<21> , \y<20> , \y<19> , \y<18> ,
         \y<17> , \y<16> , \y<15> , \y<14> , \y<13> , \y<12> , \y<11> ,
         \y<10> , \y<9> , \y<8> , \y<7> , \y<6> , \y<5> , \y<4> , \y<3> ,
         \y<2> , \y<1> , \y<0> ;
  wire   n1, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n121, n122, n123, n124, n125, n126, n127, n128,
         n129;

  OR2X2 U1 ( .A(n129), .B(\s<0> ), .Y(n121) );
  CLKINVX3 U2 ( .A(n128), .Y(n129) );
  INVX1 U3 ( .A(n128), .Y(n127) );
  INVX1 U4 ( .A(\s<1> ), .Y(n128) );
  CLKINVX3 U5 ( .A(n121), .Y(n126) );
  CLKINVX3 U6 ( .A(n124), .Y(n123) );
  CLKINVX3 U7 ( .A(n121), .Y(n125) );
  CLKINVX3 U8 ( .A(n124), .Y(n122) );
  INVX1 U9 ( .A(n3), .Y(n124) );
  NOR2BX1 U10 ( .AN(\s<0> ), .B(n129), .Y(n3) );
  OAI2BB1X1 U11 ( .A0N(\d2<1> ), .A1N(n129), .B0(n23), .Y(\y<1> ) );
  AOI22X1 U12 ( .A0(\d0<1> ), .A1(n125), .B0(\d1<1> ), .B1(n122), .Y(n23) );
  OAI2BB1X1 U13 ( .A0N(\d2<0> ), .A1N(n129), .B0(n34), .Y(\y<0> ) );
  AOI22X1 U14 ( .A0(\d0<0> ), .A1(n125), .B0(\d1<0> ), .B1(n122), .Y(n34) );
  OAI2BB1X1 U15 ( .A0N(\d2<2> ), .A1N(n129), .B0(n12), .Y(\y<2> ) );
  AOI22X1 U16 ( .A0(\d0<2> ), .A1(n126), .B0(\d1<2> ), .B1(n123), .Y(n12) );
  OAI2BB1X1 U17 ( .A0N(\d2<3> ), .A1N(n129), .B0(n9), .Y(\y<3> ) );
  AOI22X1 U18 ( .A0(\d0<3> ), .A1(n126), .B0(\d1<3> ), .B1(n123), .Y(n9) );
  OAI2BB1X1 U19 ( .A0N(\d2<4> ), .A1N(n129), .B0(n8), .Y(\y<4> ) );
  AOI22X1 U20 ( .A0(\d0<4> ), .A1(n126), .B0(\d1<4> ), .B1(n123), .Y(n8) );
  OAI2BB1X1 U21 ( .A0N(\d2<5> ), .A1N(n129), .B0(n7), .Y(\y<5> ) );
  AOI22X1 U22 ( .A0(\d0<5> ), .A1(n126), .B0(\d1<5> ), .B1(n123), .Y(n7) );
  OAI2BB1X1 U23 ( .A0N(\d2<6> ), .A1N(n129), .B0(n6), .Y(\y<6> ) );
  AOI22X1 U24 ( .A0(\d0<6> ), .A1(n126), .B0(\d1<6> ), .B1(n123), .Y(n6) );
  OAI2BB1X1 U25 ( .A0N(\d2<8> ), .A1N(n129), .B0(n4), .Y(\y<8> ) );
  AOI22X1 U26 ( .A0(\d0<8> ), .A1(n126), .B0(\d1<8> ), .B1(n123), .Y(n4) );
  OAI2BB1X1 U27 ( .A0N(\d2<10> ), .A1N(\s<1> ), .B0(n33), .Y(\y<10> ) );
  AOI22X1 U28 ( .A0(\d0<10> ), .A1(n125), .B0(\d1<10> ), .B1(n122), .Y(n33) );
  OAI2BB1X1 U29 ( .A0N(\d2<11> ), .A1N(\s<1> ), .B0(n32), .Y(\y<11> ) );
  AOI22X1 U30 ( .A0(\d0<11> ), .A1(n125), .B0(\d1<11> ), .B1(n122), .Y(n32) );
  OAI2BB1X1 U31 ( .A0N(n129), .A1N(\d2<9> ), .B0(n1), .Y(\y<9> ) );
  AOI22X1 U32 ( .A0(\d0<9> ), .A1(n126), .B0(\d1<9> ), .B1(n123), .Y(n1) );
  OAI2BB1X1 U33 ( .A0N(\d2<7> ), .A1N(n129), .B0(n5), .Y(\y<7> ) );
  AOI22X1 U34 ( .A0(\d0<7> ), .A1(n126), .B0(\d1<7> ), .B1(n123), .Y(n5) );
  OAI2BB1X1 U35 ( .A0N(\d2<15> ), .A1N(\s<1> ), .B0(n28), .Y(\y<15> ) );
  AOI22X1 U36 ( .A0(\d0<15> ), .A1(n125), .B0(\d1<15> ), .B1(n122), .Y(n28) );
  OAI2BB1X1 U37 ( .A0N(\d2<16> ), .A1N(n129), .B0(n27), .Y(\y<16> ) );
  AOI22X1 U38 ( .A0(\d0<16> ), .A1(n125), .B0(\d1<16> ), .B1(n122), .Y(n27) );
  OAI2BB1X1 U39 ( .A0N(\d2<12> ), .A1N(\s<1> ), .B0(n31), .Y(\y<12> ) );
  AOI22X1 U40 ( .A0(\d0<12> ), .A1(n125), .B0(\d1<12> ), .B1(n122), .Y(n31) );
  OAI2BB1X1 U41 ( .A0N(\d2<13> ), .A1N(\s<1> ), .B0(n30), .Y(\y<13> ) );
  AOI22X1 U42 ( .A0(\d0<13> ), .A1(n125), .B0(\d1<13> ), .B1(n122), .Y(n30) );
  OAI2BB1X1 U43 ( .A0N(\d2<14> ), .A1N(\s<1> ), .B0(n29), .Y(\y<14> ) );
  AOI22X1 U44 ( .A0(\d0<14> ), .A1(n125), .B0(\d1<14> ), .B1(n122), .Y(n29) );
  OAI2BB1X1 U45 ( .A0N(\d2<17> ), .A1N(n127), .B0(n26), .Y(\y<17> ) );
  AOI22X1 U46 ( .A0(\d0<17> ), .A1(n125), .B0(\d1<17> ), .B1(n122), .Y(n26) );
  OAI2BB1X1 U47 ( .A0N(\d2<18> ), .A1N(n127), .B0(n25), .Y(\y<18> ) );
  AOI22X1 U48 ( .A0(\d0<18> ), .A1(n125), .B0(\d1<18> ), .B1(n122), .Y(n25) );
  OAI2BB1X1 U49 ( .A0N(\d2<20> ), .A1N(n127), .B0(n22), .Y(\y<20> ) );
  AOI22X1 U50 ( .A0(\d0<20> ), .A1(n126), .B0(\d1<20> ), .B1(n123), .Y(n22) );
  OAI2BB1X1 U51 ( .A0N(\d2<22> ), .A1N(n127), .B0(n20), .Y(\y<22> ) );
  AOI22X1 U52 ( .A0(\d0<22> ), .A1(n126), .B0(\d1<22> ), .B1(n123), .Y(n20) );
  OAI2BB1X1 U53 ( .A0N(\d2<19> ), .A1N(n127), .B0(n24), .Y(\y<19> ) );
  AOI22X1 U54 ( .A0(\d0<19> ), .A1(n125), .B0(\d1<19> ), .B1(n122), .Y(n24) );
  OAI2BB1X1 U55 ( .A0N(\d2<21> ), .A1N(n127), .B0(n21), .Y(\y<21> ) );
  AOI22X1 U56 ( .A0(\d0<21> ), .A1(n126), .B0(\d1<21> ), .B1(n123), .Y(n21) );
  OAI2BB1X1 U57 ( .A0N(\d2<25> ), .A1N(n129), .B0(n17), .Y(\y<25> ) );
  AOI22X1 U58 ( .A0(\d0<25> ), .A1(n126), .B0(\d1<25> ), .B1(n123), .Y(n17) );
  OAI2BB1X1 U59 ( .A0N(\d2<24> ), .A1N(n129), .B0(n18), .Y(\y<24> ) );
  AOI22X1 U60 ( .A0(\d0<24> ), .A1(n126), .B0(\d1<24> ), .B1(n123), .Y(n18) );
  OAI2BB1X1 U61 ( .A0N(\d2<26> ), .A1N(n129), .B0(n16), .Y(\y<26> ) );
  AOI22X1 U62 ( .A0(\d0<26> ), .A1(n126), .B0(\d1<26> ), .B1(n123), .Y(n16) );
  OAI2BB1X1 U63 ( .A0N(\d2<27> ), .A1N(n129), .B0(n15), .Y(\y<27> ) );
  AOI22X1 U64 ( .A0(\d0<27> ), .A1(n126), .B0(\d1<27> ), .B1(n123), .Y(n15) );
  OAI2BB1X1 U65 ( .A0N(\d2<23> ), .A1N(n129), .B0(n19), .Y(\y<23> ) );
  AOI22X1 U66 ( .A0(\d0<23> ), .A1(n126), .B0(\d1<23> ), .B1(n123), .Y(n19) );
  OAI2BB1X1 U67 ( .A0N(\d2<28> ), .A1N(n129), .B0(n14), .Y(\y<28> ) );
  AOI22X1 U68 ( .A0(\d0<28> ), .A1(n126), .B0(\d1<28> ), .B1(n123), .Y(n14) );
  OAI2BB1X1 U69 ( .A0N(\d2<29> ), .A1N(n129), .B0(n13), .Y(\y<29> ) );
  AOI22X1 U70 ( .A0(\d0<29> ), .A1(n126), .B0(\d1<29> ), .B1(n123), .Y(n13) );
  OAI2BB1X1 U71 ( .A0N(\d2<30> ), .A1N(n129), .B0(n11), .Y(\y<30> ) );
  AOI22X1 U72 ( .A0(\d0<30> ), .A1(n126), .B0(\d1<30> ), .B1(n123), .Y(n11) );
  OAI2BB1X1 U73 ( .A0N(\d2<31> ), .A1N(n129), .B0(n10), .Y(\y<31> ) );
  AOI22X1 U74 ( .A0(\d0<31> ), .A1(n126), .B0(\d1<31> ), .B1(n123), .Y(n10) );
endmodule


module mux3_WIDTH32_1 ( .d0({\d0<31> , \d0<30> , \d0<29> , \d0<28> , \d0<27> , 
        \d0<26> , \d0<25> , \d0<24> , \d0<23> , \d0<22> , \d0<21> , \d0<20> , 
        \d0<19> , \d0<18> , \d0<17> , \d0<16> , \d0<15> , \d0<14> , \d0<13> , 
        \d0<12> , \d0<11> , \d0<10> , \d0<9> , \d0<8> , \d0<7> , \d0<6> , 
        \d0<5> , \d0<4> , \d0<3> , \d0<2> , \d0<1> , \d0<0> }), .d1({\d1<31> , 
        \d1<30> , \d1<29> , \d1<28> , \d1<27> , \d1<26> , \d1<25> , \d1<24> , 
        \d1<23> , \d1<22> , \d1<21> , \d1<20> , \d1<19> , \d1<18> , \d1<17> , 
        \d1<16> , \d1<15> , \d1<14> , \d1<13> , \d1<12> , \d1<11> , \d1<10> , 
        \d1<9> , \d1<8> , \d1<7> , \d1<6> , \d1<5> , \d1<4> , \d1<3> , \d1<2> , 
        \d1<1> , \d1<0> }), .d2({\d2<31> , \d2<30> , \d2<29> , \d2<28> , 
        \d2<27> , \d2<26> , \d2<25> , \d2<24> , \d2<23> , \d2<22> , \d2<21> , 
        \d2<20> , \d2<19> , \d2<18> , \d2<17> , \d2<16> , \d2<15> , \d2<14> , 
        \d2<13> , \d2<12> , \d2<11> , \d2<10> , \d2<9> , \d2<8> , \d2<7> , 
        \d2<6> , \d2<5> , \d2<4> , \d2<3> , \d2<2> , \d2<1> , \d2<0> }), .s({
        \s<1> , \s<0> }), .y({\y<31> , \y<30> , \y<29> , \y<28> , \y<27> , 
        \y<26> , \y<25> , \y<24> , \y<23> , \y<22> , \y<21> , \y<20> , \y<19> , 
        \y<18> , \y<17> , \y<16> , \y<15> , \y<14> , \y<13> , \y<12> , \y<11> , 
        \y<10> , \y<9> , \y<8> , \y<7> , \y<6> , \y<5> , \y<4> , \y<3> , 
        \y<2> , \y<1> , \y<0> }) );
  input \d0<31> , \d0<30> , \d0<29> , \d0<28> , \d0<27> , \d0<26> , \d0<25> ,
         \d0<24> , \d0<23> , \d0<22> , \d0<21> , \d0<20> , \d0<19> , \d0<18> ,
         \d0<17> , \d0<16> , \d0<15> , \d0<14> , \d0<13> , \d0<12> , \d0<11> ,
         \d0<10> , \d0<9> , \d0<8> , \d0<7> , \d0<6> , \d0<5> , \d0<4> ,
         \d0<3> , \d0<2> , \d0<1> , \d0<0> , \d1<31> , \d1<30> , \d1<29> ,
         \d1<28> , \d1<27> , \d1<26> , \d1<25> , \d1<24> , \d1<23> , \d1<22> ,
         \d1<21> , \d1<20> , \d1<19> , \d1<18> , \d1<17> , \d1<16> , \d1<15> ,
         \d1<14> , \d1<13> , \d1<12> , \d1<11> , \d1<10> , \d1<9> , \d1<8> ,
         \d1<7> , \d1<6> , \d1<5> , \d1<4> , \d1<3> , \d1<2> , \d1<1> ,
         \d1<0> , \d2<31> , \d2<30> , \d2<29> , \d2<28> , \d2<27> , \d2<26> ,
         \d2<25> , \d2<24> , \d2<23> , \d2<22> , \d2<21> , \d2<20> , \d2<19> ,
         \d2<18> , \d2<17> , \d2<16> , \d2<15> , \d2<14> , \d2<13> , \d2<12> ,
         \d2<11> , \d2<10> , \d2<9> , \d2<8> , \d2<7> , \d2<6> , \d2<5> ,
         \d2<4> , \d2<3> , \d2<2> , \d2<1> , \d2<0> , \s<1> , \s<0> ;
  output \y<31> , \y<30> , \y<29> , \y<28> , \y<27> , \y<26> , \y<25> ,
         \y<24> , \y<23> , \y<22> , \y<21> , \y<20> , \y<19> , \y<18> ,
         \y<17> , \y<16> , \y<15> , \y<14> , \y<13> , \y<12> , \y<11> ,
         \y<10> , \y<9> , \y<8> , \y<7> , \y<6> , \y<5> , \y<4> , \y<3> ,
         \y<2> , \y<1> , \y<0> ;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n121, n122, n123, n124, n125, n126, n127, n128,
         n129;

  CLKINVX3 U1 ( .A(n128), .Y(n129) );
  INVX1 U2 ( .A(n128), .Y(n127) );
  INVX1 U3 ( .A(\s<1> ), .Y(n128) );
  CLKINVX3 U4 ( .A(n126), .Y(n124) );
  CLKINVX3 U5 ( .A(n123), .Y(n121) );
  CLKINVX3 U6 ( .A(n126), .Y(n125) );
  CLKINVX3 U7 ( .A(n123), .Y(n122) );
  INVX1 U8 ( .A(n3), .Y(n123) );
  INVX1 U9 ( .A(n2), .Y(n126) );
  NOR2X1 U10 ( .A(n129), .B(\s<0> ), .Y(n2) );
  NOR2BX1 U11 ( .AN(\s<0> ), .B(n129), .Y(n3) );
  OAI2BB1X1 U12 ( .A0N(\d2<31> ), .A1N(n129), .B0(n10), .Y(\y<31> ) );
  AOI22X1 U13 ( .A0(\d0<31> ), .A1(n125), .B0(\d1<31> ), .B1(n122), .Y(n10) );
  OAI2BB1X1 U14 ( .A0N(\d2<26> ), .A1N(\s<1> ), .B0(n16), .Y(\y<26> ) );
  AOI22X1 U15 ( .A0(\d0<26> ), .A1(n124), .B0(\d1<26> ), .B1(n121), .Y(n16) );
  OAI2BB1X1 U16 ( .A0N(\d2<27> ), .A1N(n129), .B0(n15), .Y(\y<27> ) );
  AOI22X1 U17 ( .A0(\d0<27> ), .A1(n124), .B0(\d1<27> ), .B1(n121), .Y(n15) );
  OAI2BB1X1 U18 ( .A0N(\d2<28> ), .A1N(n129), .B0(n14), .Y(\y<28> ) );
  AOI22X1 U19 ( .A0(\d0<28> ), .A1(n124), .B0(\d1<28> ), .B1(n121), .Y(n14) );
  OAI2BB1X1 U20 ( .A0N(\d2<29> ), .A1N(n129), .B0(n13), .Y(\y<29> ) );
  AOI22X1 U21 ( .A0(\d0<29> ), .A1(n124), .B0(\d1<29> ), .B1(n121), .Y(n13) );
  OAI2BB1X1 U22 ( .A0N(\d2<30> ), .A1N(n129), .B0(n11), .Y(\y<30> ) );
  AOI22X1 U23 ( .A0(\d0<30> ), .A1(n124), .B0(\d1<30> ), .B1(n121), .Y(n11) );
  OAI2BB1X1 U24 ( .A0N(\d2<21> ), .A1N(n127), .B0(n21), .Y(\y<21> ) );
  AOI22X1 U25 ( .A0(\d0<21> ), .A1(n124), .B0(\d1<21> ), .B1(n121), .Y(n21) );
  OAI2BB1X1 U26 ( .A0N(\d2<22> ), .A1N(n129), .B0(n20), .Y(\y<22> ) );
  AOI22X1 U27 ( .A0(\d0<22> ), .A1(n124), .B0(\d1<22> ), .B1(n121), .Y(n20) );
  OAI2BB1X1 U28 ( .A0N(\d2<23> ), .A1N(n129), .B0(n19), .Y(\y<23> ) );
  AOI22X1 U29 ( .A0(\d0<23> ), .A1(n124), .B0(\d1<23> ), .B1(n121), .Y(n19) );
  OAI2BB1X1 U30 ( .A0N(\d2<24> ), .A1N(n129), .B0(n18), .Y(\y<24> ) );
  AOI22X1 U31 ( .A0(\d0<24> ), .A1(n124), .B0(\d1<24> ), .B1(n121), .Y(n18) );
  OAI2BB1X1 U32 ( .A0N(\d2<25> ), .A1N(\s<1> ), .B0(n17), .Y(\y<25> ) );
  AOI22X1 U33 ( .A0(\d0<25> ), .A1(n124), .B0(\d1<25> ), .B1(n121), .Y(n17) );
  OAI2BB1X1 U34 ( .A0N(\d2<17> ), .A1N(\s<1> ), .B0(n26), .Y(\y<17> ) );
  AOI22X1 U35 ( .A0(\d0<17> ), .A1(n125), .B0(\d1<17> ), .B1(n122), .Y(n26) );
  OAI2BB1X1 U36 ( .A0N(\d2<18> ), .A1N(n129), .B0(n25), .Y(\y<18> ) );
  AOI22X1 U37 ( .A0(\d0<18> ), .A1(n124), .B0(\d1<18> ), .B1(n121), .Y(n25) );
  OAI2BB1X1 U38 ( .A0N(\d2<19> ), .A1N(n127), .B0(n24), .Y(\y<19> ) );
  AOI22X1 U39 ( .A0(\d0<19> ), .A1(n124), .B0(\d1<19> ), .B1(n121), .Y(n24) );
  OAI2BB1X1 U40 ( .A0N(\d2<20> ), .A1N(\s<1> ), .B0(n22), .Y(\y<20> ) );
  AOI22X1 U41 ( .A0(\d0<20> ), .A1(n124), .B0(\d1<20> ), .B1(n121), .Y(n22) );
  OAI2BB1X1 U42 ( .A0N(\d2<12> ), .A1N(n127), .B0(n31), .Y(\y<12> ) );
  AOI22X1 U43 ( .A0(\d0<12> ), .A1(n125), .B0(\d1<12> ), .B1(n122), .Y(n31) );
  OAI2BB1X1 U44 ( .A0N(\d2<13> ), .A1N(n127), .B0(n30), .Y(\y<13> ) );
  AOI22X1 U45 ( .A0(\d0<13> ), .A1(n124), .B0(\d1<13> ), .B1(n121), .Y(n30) );
  OAI2BB1X1 U46 ( .A0N(\d2<14> ), .A1N(n127), .B0(n29), .Y(\y<14> ) );
  AOI22X1 U47 ( .A0(\d0<14> ), .A1(n125), .B0(\d1<14> ), .B1(n121), .Y(n29) );
  OAI2BB1X1 U48 ( .A0N(\d2<15> ), .A1N(n129), .B0(n28), .Y(\y<15> ) );
  AOI22X1 U49 ( .A0(\d0<15> ), .A1(n124), .B0(\d1<15> ), .B1(n121), .Y(n28) );
  OAI2BB1X1 U50 ( .A0N(\d2<16> ), .A1N(n127), .B0(n27), .Y(\y<16> ) );
  AOI22X1 U51 ( .A0(\d0<16> ), .A1(n124), .B0(\d1<16> ), .B1(n121), .Y(n27) );
  OAI2BB1X1 U52 ( .A0N(n129), .A1N(\d2<9> ), .B0(n1), .Y(\y<9> ) );
  AOI22X1 U53 ( .A0(\d0<9> ), .A1(n125), .B0(\d1<9> ), .B1(n122), .Y(n1) );
  OAI2BB1X1 U54 ( .A0N(\d2<7> ), .A1N(n129), .B0(n5), .Y(\y<7> ) );
  AOI22X1 U55 ( .A0(\d0<7> ), .A1(n125), .B0(\d1<7> ), .B1(n122), .Y(n5) );
  OAI2BB1X1 U56 ( .A0N(\d2<8> ), .A1N(n129), .B0(n4), .Y(\y<8> ) );
  AOI22X1 U57 ( .A0(\d0<8> ), .A1(n125), .B0(\d1<8> ), .B1(n122), .Y(n4) );
  OAI2BB1X1 U58 ( .A0N(\d2<10> ), .A1N(\s<1> ), .B0(n33), .Y(\y<10> ) );
  AOI22X1 U59 ( .A0(\d0<10> ), .A1(n124), .B0(\d1<10> ), .B1(n121), .Y(n33) );
  OAI2BB1X1 U60 ( .A0N(\d2<11> ), .A1N(\s<1> ), .B0(n32), .Y(\y<11> ) );
  AOI22X1 U61 ( .A0(\d0<11> ), .A1(n125), .B0(\d1<11> ), .B1(n122), .Y(n32) );
  OAI2BB1X1 U62 ( .A0N(\d2<2> ), .A1N(n129), .B0(n12), .Y(\y<2> ) );
  AOI22X1 U63 ( .A0(\d0<2> ), .A1(n124), .B0(\d1<2> ), .B1(n121), .Y(n12) );
  OAI2BB1X1 U64 ( .A0N(\d2<3> ), .A1N(n129), .B0(n9), .Y(\y<3> ) );
  AOI22X1 U65 ( .A0(\d0<3> ), .A1(n125), .B0(\d1<3> ), .B1(n122), .Y(n9) );
  OAI2BB1X1 U66 ( .A0N(\d2<4> ), .A1N(n129), .B0(n8), .Y(\y<4> ) );
  AOI22X1 U67 ( .A0(\d0<4> ), .A1(n125), .B0(\d1<4> ), .B1(n122), .Y(n8) );
  OAI2BB1X1 U68 ( .A0N(\d2<5> ), .A1N(n129), .B0(n7), .Y(\y<5> ) );
  AOI22X1 U69 ( .A0(\d0<5> ), .A1(n125), .B0(\d1<5> ), .B1(n122), .Y(n7) );
  OAI2BB1X1 U70 ( .A0N(\d2<6> ), .A1N(n129), .B0(n6), .Y(\y<6> ) );
  AOI22X1 U71 ( .A0(\d0<6> ), .A1(n125), .B0(\d1<6> ), .B1(n122), .Y(n6) );
  OAI2BB1X1 U72 ( .A0N(\d2<1> ), .A1N(n129), .B0(n23), .Y(\y<1> ) );
  AOI22X1 U73 ( .A0(\d0<1> ), .A1(n124), .B0(\d1<1> ), .B1(n122), .Y(n23) );
  OAI2BB1X1 U74 ( .A0N(\d2<0> ), .A1N(n129), .B0(n34), .Y(\y<0> ) );
  AOI22X1 U75 ( .A0(\d0<0> ), .A1(n2), .B0(\d1<0> ), .B1(n121), .Y(n34) );
endmodule


module regfile ( clk, we3, .ra1({\ra1<3> , \ra1<2> , \ra1<1> , \ra1<0> }), 
    .ra2({\ra2<3> , \ra2<2> , \ra2<1> , \ra2<0> }), .wa3({\wa3<3> , \wa3<2> , 
        \wa3<1> , \wa3<0> }), .wd3({\wd3<31> , \wd3<30> , \wd3<29> , \wd3<28> , 
        \wd3<27> , \wd3<26> , \wd3<25> , \wd3<24> , \wd3<23> , \wd3<22> , 
        \wd3<21> , \wd3<20> , \wd3<19> , \wd3<18> , \wd3<17> , \wd3<16> , 
        \wd3<15> , \wd3<14> , \wd3<13> , \wd3<12> , \wd3<11> , \wd3<10> , 
        \wd3<9> , \wd3<8> , \wd3<7> , \wd3<6> , \wd3<5> , \wd3<4> , \wd3<3> , 
        \wd3<2> , \wd3<1> , \wd3<0> }), .r15({\r15<31> , \r15<30> , \r15<29> , 
        \r15<28> , \r15<27> , \r15<26> , \r15<25> , \r15<24> , \r15<23> , 
        \r15<22> , \r15<21> , \r15<20> , \r15<19> , \r15<18> , \r15<17> , 
        \r15<16> , \r15<15> , \r15<14> , \r15<13> , \r15<12> , \r15<11> , 
        \r15<10> , \r15<9> , \r15<8> , \r15<7> , \r15<6> , \r15<5> , \r15<4> , 
        \r15<3> , \r15<2> , \r15<1> , \r15<0> }), .rd1({\rd1<31> , \rd1<30> , 
        \rd1<29> , \rd1<28> , \rd1<27> , \rd1<26> , \rd1<25> , \rd1<24> , 
        \rd1<23> , \rd1<22> , \rd1<21> , \rd1<20> , \rd1<19> , \rd1<18> , 
        \rd1<17> , \rd1<16> , \rd1<15> , \rd1<14> , \rd1<13> , \rd1<12> , 
        \rd1<11> , \rd1<10> , \rd1<9> , \rd1<8> , \rd1<7> , \rd1<6> , \rd1<5> , 
        \rd1<4> , \rd1<3> , \rd1<2> , \rd1<1> , \rd1<0> }), .rd2({\rd2<31> , 
        \rd2<30> , \rd2<29> , \rd2<28> , \rd2<27> , \rd2<26> , \rd2<25> , 
        \rd2<24> , \rd2<23> , \rd2<22> , \rd2<21> , \rd2<20> , \rd2<19> , 
        \rd2<18> , \rd2<17> , \rd2<16> , \rd2<15> , \rd2<14> , \rd2<13> , 
        \rd2<12> , \rd2<11> , \rd2<10> , \rd2<9> , \rd2<8> , \rd2<7> , 
        \rd2<6> , \rd2<5> , \rd2<4> , \rd2<3> , \rd2<2> , \rd2<1> , \rd2<0> })
 );
  input clk, we3, \ra1<3> , \ra1<2> , \ra1<1> , \ra1<0> , \ra2<3> , \ra2<2> ,
         \ra2<1> , \ra2<0> , \wa3<3> , \wa3<2> , \wa3<1> , \wa3<0> , \wd3<31> ,
         \wd3<30> , \wd3<29> , \wd3<28> , \wd3<27> , \wd3<26> , \wd3<25> ,
         \wd3<24> , \wd3<23> , \wd3<22> , \wd3<21> , \wd3<20> , \wd3<19> ,
         \wd3<18> , \wd3<17> , \wd3<16> , \wd3<15> , \wd3<14> , \wd3<13> ,
         \wd3<12> , \wd3<11> , \wd3<10> , \wd3<9> , \wd3<8> , \wd3<7> ,
         \wd3<6> , \wd3<5> , \wd3<4> , \wd3<3> , \wd3<2> , \wd3<1> , \wd3<0> ,
         \r15<31> , \r15<30> , \r15<29> , \r15<28> , \r15<27> , \r15<26> ,
         \r15<25> , \r15<24> , \r15<23> , \r15<22> , \r15<21> , \r15<20> ,
         \r15<19> , \r15<18> , \r15<17> , \r15<16> , \r15<15> , \r15<14> ,
         \r15<13> , \r15<12> , \r15<11> , \r15<10> , \r15<9> , \r15<8> ,
         \r15<7> , \r15<6> , \r15<5> , \r15<4> , \r15<3> , \r15<2> , \r15<1> ,
         \r15<0> ;
  output \rd1<31> , \rd1<30> , \rd1<29> , \rd1<28> , \rd1<27> , \rd1<26> ,
         \rd1<25> , \rd1<24> , \rd1<23> , \rd1<22> , \rd1<21> , \rd1<20> ,
         \rd1<19> , \rd1<18> , \rd1<17> , \rd1<16> , \rd1<15> , \rd1<14> ,
         \rd1<13> , \rd1<12> , \rd1<11> , \rd1<10> , \rd1<9> , \rd1<8> ,
         \rd1<7> , \rd1<6> , \rd1<5> , \rd1<4> , \rd1<3> , \rd1<2> , \rd1<1> ,
         \rd1<0> , \rd2<31> , \rd2<30> , \rd2<29> , \rd2<28> , \rd2<27> ,
         \rd2<26> , \rd2<25> , \rd2<24> , \rd2<23> , \rd2<22> , \rd2<21> ,
         \rd2<20> , \rd2<19> , \rd2<18> , \rd2<17> , \rd2<16> , \rd2<15> ,
         \rd2<14> , \rd2<13> , \rd2<12> , \rd2<11> , \rd2<10> , \rd2<9> ,
         \rd2<8> , \rd2<7> , \rd2<6> , \rd2<5> , \rd2<4> , \rd2<3> , \rd2<2> ,
         \rd2<1> , \rd2<0> ;
  wire   N12, N13, N14, N15, N16, N17, N18, N19, \rf<11><31> , \rf<11><30> ,
         \rf<11><29> , \rf<11><28> , \rf<11><27> , \rf<11><26> , \rf<11><25> ,
         \rf<11><24> , \rf<11><23> , \rf<11><22> , \rf<11><21> , \rf<11><20> ,
         \rf<11><19> , \rf<11><18> , \rf<11><17> , \rf<11><16> , \rf<11><15> ,
         \rf<11><14> , \rf<11><13> , \rf<11><12> , \rf<11><11> , \rf<11><10> ,
         \rf<11><9> , \rf<11><8> , \rf<11><7> , \rf<11><6> , \rf<11><5> ,
         \rf<11><4> , \rf<11><3> , \rf<11><2> , \rf<11><1> , \rf<11><0> ,
         \rf<10><31> , \rf<10><30> , \rf<10><29> , \rf<10><28> , \rf<10><27> ,
         \rf<10><26> , \rf<10><25> , \rf<10><24> , \rf<10><23> , \rf<10><22> ,
         \rf<10><21> , \rf<10><20> , \rf<10><19> , \rf<10><18> , \rf<10><17> ,
         \rf<10><16> , \rf<10><15> , \rf<10><14> , \rf<10><13> , \rf<10><12> ,
         \rf<10><11> , \rf<10><10> , \rf<10><9> , \rf<10><8> , \rf<10><7> ,
         \rf<10><6> , \rf<10><5> , \rf<10><4> , \rf<10><3> , \rf<10><2> ,
         \rf<10><1> , \rf<10><0> , \rf<7><31> , \rf<7><30> , \rf<7><29> ,
         \rf<7><28> , \rf<7><27> , \rf<7><26> , \rf<7><25> , \rf<7><24> ,
         \rf<7><23> , \rf<7><22> , \rf<7><21> , \rf<7><20> , \rf<7><19> ,
         \rf<7><18> , \rf<7><17> , \rf<7><16> , \rf<7><15> , \rf<7><14> ,
         \rf<7><13> , \rf<7><12> , \rf<7><11> , \rf<7><10> , \rf<7><9> ,
         \rf<7><8> , \rf<7><7> , \rf<7><6> , \rf<7><5> , \rf<7><4> ,
         \rf<7><3> , \rf<7><2> , \rf<7><1> , \rf<7><0> , \rf<6><31> ,
         \rf<6><30> , \rf<6><29> , \rf<6><28> , \rf<6><27> , \rf<6><26> ,
         \rf<6><25> , \rf<6><24> , \rf<6><23> , \rf<6><22> , \rf<6><21> ,
         \rf<6><20> , \rf<6><19> , \rf<6><18> , \rf<6><17> , \rf<6><16> ,
         \rf<6><15> , \rf<6><14> , \rf<6><13> , \rf<6><12> , \rf<6><11> ,
         \rf<6><10> , \rf<6><9> , \rf<6><8> , \rf<6><7> , \rf<6><6> ,
         \rf<6><5> , \rf<6><4> , \rf<6><3> , \rf<6><2> , \rf<6><1> ,
         \rf<6><0> , \rf<2><31> , \rf<2><30> , \rf<2><29> , \rf<2><28> ,
         \rf<2><27> , \rf<2><26> , \rf<2><25> , \rf<2><24> , \rf<2><23> ,
         \rf<2><22> , \rf<2><21> , \rf<2><20> , \rf<2><19> , \rf<2><18> ,
         \rf<2><17> , \rf<2><16> , \rf<2><15> , \rf<2><14> , \rf<2><13> ,
         \rf<2><12> , \rf<2><11> , \rf<2><10> , \rf<2><9> , \rf<2><8> ,
         \rf<2><7> , \rf<2><6> , \rf<2><5> , \rf<2><4> , \rf<2><3> ,
         \rf<2><2> , \rf<2><1> , \rf<2><0> , n13, n15, n16, n1579, n1580,
         n3939, n3940, n3941, n3942, n3943, n3944, n3945, n3946, n3947, n3948,
         n3949, n3950, n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3958,
         n3959, n3960, n3961, n3962, n3963, n3964, n3965, n3966, n3967, n3968,
         n3969, n3970, n3971, n3972, n3973, n3974, n3975, n3976, n3977, n3978,
         n3979, n3980, n3981, n3982, n3983, n3984, n3985, n3986, n3987, n3988,
         n3989, n3990, n3991, n3992, n3993, n3994, n3995, n3996, n3997, n3998,
         n3999, n4000, n4001, n4002, n4003, n4004, n4005, n4006, n4007, n4008,
         n4009, n4010, n4011, n4012, n4013, n4014, n4015, n4016, n4017, n4018,
         n4019, n4020, n4021, n4022, n4023, n4024, n4025, n4026, n4027, n4028,
         n4029, n4030, n4031, n4032, n4033, n4034, n4099, n4100, n4101, n4102,
         n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112,
         n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122,
         n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132,
         n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142,
         n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152,
         n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162,
         n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172,
         n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182,
         n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192,
         n4193, n4194, n4291, n4292, n4293, n4294, n4295, n4296, n4297, n4298,
         n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4306, n4307, n4308,
         n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4318,
         n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328,
         n4329, n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337, n4338,
         n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4348,
         n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358,
         n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368,
         n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378,
         n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388,
         n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398,
         n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408,
         n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418,
         n1008, n1009, n1010, n1011, n1014, n1019, n1024, n1028, n1029, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
         n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
         n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
         n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
         n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
         n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
         n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
         n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
         n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
         n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
         n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
         n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
         n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
         n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
         n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
         n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
         n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
         n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
         n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
         n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
         n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
         n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
         n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
         n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
         n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
         n1283, n1284, n1285, n1286, n1287, n1290, n1291, n1292, n1295, n1296,
         n1297, n1300, n1301, n1302, n1304, n1305, n1306, n1307, n1308, n1309,
         n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319,
         n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329,
         n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339,
         n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349,
         n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359,
         n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369,
         n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379,
         n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389,
         n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399,
         n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409,
         n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419,
         n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429,
         n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439,
         n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449,
         n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459,
         n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469,
         n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479,
         n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489,
         n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499,
         n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509,
         n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519,
         n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529,
         n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539,
         n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549,
         n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559,
         n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569,
         n1570, n1571, n1572, n1573, n1574, n1575, n4602, n4603, n4604, n4605,
         n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615,
         n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624, n4625,
         n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634, n4635,
         n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644, n4645,
         n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654, n4655,
         n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664, n4665,
         n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674, n4675,
         n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685,
         n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694, n4695,
         n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705,
         n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714, n4715,
         n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724, n4725,
         n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734, n4735,
         n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744, n4745,
         n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755,
         n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4765,
         n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774, n4775,
         n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784, n4785,
         n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794, n4795,
         n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804, n4805,
         n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814, n4815,
         n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824, n4825,
         n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4835,
         n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844, n4845,
         n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854, n4855,
         n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864, n4865,
         n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4875,
         n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885,
         n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894, n4895,
         n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904, n4905,
         n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914, n4915,
         n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924, n4925,
         n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934, n4935,
         n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944, n4945,
         n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954, n4955,
         n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964, n4965,
         n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974, n4975,
         n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984, n4985,
         n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994, n4995,
         n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004, n5005,
         n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014, n5015,
         n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024, n5025,
         n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034, n5035,
         n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044, n5045,
         n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054, n5055,
         n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064, n5065,
         n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074, n5075,
         n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084, n5085,
         n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094, n5095,
         n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103, n5104, n5105,
         n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114, n5115,
         n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123, n5124, n5125,
         n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134, n5135,
         n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143, n5144, n5145,
         n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153, n5154, n5155,
         n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163, n5164, n5165,
         n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173, n5174, n5175,
         n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183, n5184, n5185,
         n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193, n5194, n5195,
         n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203, n5204, n5205,
         n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213, n5214, n5215,
         n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223, n5224, n5225,
         n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233, n5234, n5235,
         n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243, n5244, n5245,
         n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253, n5254, n5255,
         n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263, n5264, n5265,
         n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273, n5274, n5275,
         n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283, n5284, n5285,
         n5286, n5287, n5288, n5289, n5290;
  assign N12 = \ra1<0> ;
  assign N13 = \ra1<1> ;
  assign N14 = \ra1<2> ;
  assign N15 = \ra1<3> ;
  assign N16 = \ra2<0> ;
  assign N17 = \ra2<1> ;
  assign N18 = \ra2<2> ;
  assign N19 = \ra2<3> ;

  EDFFX1 \rf_reg<4><31>  ( .D(n5141), .E(n5146), .CK(clk), .Q(n4980), .QN(
        n3940) );
  EDFFX1 \rf_reg<4><30>  ( .D(n5140), .E(n5146), .CK(clk), .Q(n4977), .QN(
        n3943) );
  EDFFX1 \rf_reg<4><29>  ( .D(n5139), .E(n5146), .CK(clk), .Q(n4974), .QN(
        n3958) );
  EDFFX1 \rf_reg<4><28>  ( .D(n5138), .E(n5146), .CK(clk), .Q(n4971), .QN(
        n3956) );
  EDFFX1 \rf_reg<4><27>  ( .D(n5137), .E(n5146), .CK(clk), .Q(n4968), .QN(
        n3954) );
  EDFFX1 \rf_reg<4><26>  ( .D(n5136), .E(n5146), .CK(clk), .Q(n4965), .QN(
        n3952) );
  EDFFX1 \rf_reg<4><25>  ( .D(n5135), .E(n5146), .CK(clk), .Q(n4962), .QN(
        n3950) );
  EDFFX1 \rf_reg<4><24>  ( .D(n5134), .E(n5146), .CK(clk), .Q(n4959), .QN(
        n3973) );
  EDFFX1 \rf_reg<4><23>  ( .D(n5133), .E(n5146), .CK(clk), .Q(n4956), .QN(
        n3971) );
  EDFFX1 \rf_reg<4><22>  ( .D(n5132), .E(n5146), .CK(clk), .Q(n4953), .QN(
        n3969) );
  EDFFX1 \rf_reg<4><21>  ( .D(n5131), .E(n5146), .CK(clk), .Q(n4950), .QN(
        n3967) );
  EDFFX1 \rf_reg<4><20>  ( .D(n5130), .E(n5146), .CK(clk), .Q(n4947), .QN(
        n3965) );
  EDFFX1 \rf_reg<4><19>  ( .D(n5129), .E(n5147), .CK(clk), .Q(n4944), .QN(
        n3988) );
  EDFFX1 \rf_reg<4><18>  ( .D(n5128), .E(n5147), .CK(clk), .Q(n4941), .QN(
        n3986) );
  EDFFX1 \rf_reg<4><17>  ( .D(n5127), .E(n5147), .CK(clk), .Q(n4938), .QN(
        n3984) );
  EDFFX1 \rf_reg<4><16>  ( .D(n5126), .E(n5147), .CK(clk), .Q(n4935), .QN(
        n3982) );
  EDFFX1 \rf_reg<4><15>  ( .D(n5125), .E(n5147), .CK(clk), .Q(n4932), .QN(
        n3980) );
  EDFFX1 \rf_reg<4><14>  ( .D(n5124), .E(n5147), .CK(clk), .Q(n4929), .QN(
        n4006) );
  EDFFX1 \rf_reg<4><13>  ( .D(n5123), .E(n5147), .CK(clk), .Q(n4926), .QN(
        n4004) );
  EDFFX1 \rf_reg<4><12>  ( .D(n5122), .E(n5147), .CK(clk), .Q(n4923), .QN(
        n4002) );
  EDFFX1 \rf_reg<4><11>  ( .D(n5121), .E(n5147), .CK(clk), .Q(n4920), .QN(
        n4000) );
  EDFFX1 \rf_reg<4><10>  ( .D(n5120), .E(n5147), .CK(clk), .Q(n4917), .QN(
        n3998) );
  EDFFX1 \rf_reg<4><9>  ( .D(n5119), .E(n5147), .CK(clk), .Q(n4914), .QN(n3996) );
  EDFFX1 \rf_reg<4><8>  ( .D(n5118), .E(n5147), .CK(clk), .Q(n4911), .QN(n4021) );
  EDFFX1 \rf_reg<4><7>  ( .D(n5117), .E(n1574), .CK(clk), .Q(n4908), .QN(n4019) );
  EDFFX1 \rf_reg<4><6>  ( .D(n5116), .E(n1574), .CK(clk), .Q(n4905), .QN(n4017) );
  EDFFX1 \rf_reg<4><5>  ( .D(n5115), .E(n5146), .CK(clk), .Q(n4902), .QN(n4015) );
  EDFFX1 \rf_reg<4><4>  ( .D(n5114), .E(n5147), .CK(clk), .Q(n4899), .QN(n4013) );
  EDFFX1 \rf_reg<4><3>  ( .D(n5113), .E(n5146), .CK(clk), .Q(n4896), .QN(n4033) );
  EDFFX1 \rf_reg<4><2>  ( .D(n5112), .E(n5147), .CK(clk), .Q(n4893), .QN(n4031) );
  EDFFX1 \rf_reg<4><1>  ( .D(n5111), .E(n5146), .CK(clk), .Q(n4890), .QN(n4029) );
  EDFFX1 \rf_reg<4><0>  ( .D(n5110), .E(n5147), .CK(clk), .Q(n4887), .QN(n4027) );
  EDFFX1 \rf_reg<12><31>  ( .D(n5141), .E(n5230), .CK(clk), .Q(n4979), .QN(
        n4322) );
  EDFFX1 \rf_reg<12><30>  ( .D(n5140), .E(n5230), .CK(clk), .Q(n4976), .QN(
        n4321) );
  EDFFX1 \rf_reg<12><29>  ( .D(n5139), .E(n5230), .CK(clk), .Q(n4973), .QN(
        n4320) );
  EDFFX1 \rf_reg<12><28>  ( .D(n5138), .E(n5230), .CK(clk), .Q(n4970), .QN(
        n4319) );
  EDFFX1 \rf_reg<12><27>  ( .D(n5137), .E(n5230), .CK(clk), .Q(n4967), .QN(
        n4318) );
  EDFFX1 \rf_reg<12><26>  ( .D(n5136), .E(n5230), .CK(clk), .Q(n4964), .QN(
        n4317) );
  EDFFX1 \rf_reg<12><25>  ( .D(n5135), .E(n5230), .CK(clk), .Q(n4961), .QN(
        n4316) );
  EDFFX1 \rf_reg<12><24>  ( .D(n5134), .E(n5230), .CK(clk), .Q(n4958), .QN(
        n4315) );
  EDFFX1 \rf_reg<12><23>  ( .D(n5133), .E(n5230), .CK(clk), .Q(n4955), .QN(
        n4314) );
  EDFFX1 \rf_reg<12><22>  ( .D(n5132), .E(n5230), .CK(clk), .Q(n4952), .QN(
        n4313) );
  EDFFX1 \rf_reg<12><21>  ( .D(n5131), .E(n5230), .CK(clk), .Q(n4949), .QN(
        n4312) );
  EDFFX1 \rf_reg<12><20>  ( .D(n5130), .E(n5230), .CK(clk), .Q(n4946), .QN(
        n4311) );
  EDFFX1 \rf_reg<12><19>  ( .D(n5129), .E(n5231), .CK(clk), .Q(n4943), .QN(
        n4310) );
  EDFFX1 \rf_reg<12><18>  ( .D(n5128), .E(n5231), .CK(clk), .Q(n4940), .QN(
        n4309) );
  EDFFX1 \rf_reg<12><17>  ( .D(n5127), .E(n5231), .CK(clk), .Q(n4937), .QN(
        n4308) );
  EDFFX1 \rf_reg<12><16>  ( .D(n5126), .E(n5231), .CK(clk), .Q(n4934), .QN(
        n4307) );
  EDFFX1 \rf_reg<12><15>  ( .D(n5125), .E(n5231), .CK(clk), .Q(n4931), .QN(
        n4306) );
  EDFFX1 \rf_reg<12><14>  ( .D(n5124), .E(n5231), .CK(clk), .Q(n4928), .QN(
        n4305) );
  EDFFX1 \rf_reg<12><13>  ( .D(n5123), .E(n5231), .CK(clk), .Q(n4925), .QN(
        n4304) );
  EDFFX1 \rf_reg<12><12>  ( .D(n5122), .E(n5231), .CK(clk), .Q(n4922), .QN(
        n4303) );
  EDFFX1 \rf_reg<12><11>  ( .D(n5121), .E(n5231), .CK(clk), .Q(n4919), .QN(
        n4302) );
  EDFFX1 \rf_reg<12><10>  ( .D(n5120), .E(n5231), .CK(clk), .Q(n4916), .QN(
        n4301) );
  EDFFX1 \rf_reg<12><9>  ( .D(n5119), .E(n5231), .CK(clk), .Q(n4913), .QN(
        n4300) );
  EDFFX1 \rf_reg<12><8>  ( .D(n5118), .E(n5231), .CK(clk), .Q(n4910), .QN(
        n4299) );
  EDFFX1 \rf_reg<12><7>  ( .D(n5117), .E(n1579), .CK(clk), .Q(n4907), .QN(
        n4298) );
  EDFFX1 \rf_reg<12><6>  ( .D(n5116), .E(n1579), .CK(clk), .Q(n4904), .QN(
        n4297) );
  EDFFX1 \rf_reg<12><5>  ( .D(n5115), .E(n5230), .CK(clk), .Q(n4901), .QN(
        n4296) );
  EDFFX1 \rf_reg<12><4>  ( .D(n5114), .E(n5231), .CK(clk), .Q(n4898), .QN(
        n4295) );
  EDFFX1 \rf_reg<12><3>  ( .D(n5113), .E(n5230), .CK(clk), .Q(n4895), .QN(
        n4294) );
  EDFFX1 \rf_reg<12><2>  ( .D(n5112), .E(n5231), .CK(clk), .Q(n4892), .QN(
        n4293) );
  EDFFX1 \rf_reg<12><1>  ( .D(n5111), .E(n5230), .CK(clk), .Q(n4889), .QN(
        n4292) );
  EDFFX1 \rf_reg<12><0>  ( .D(n5110), .E(n5231), .CK(clk), .Q(n4886), .QN(
        n4291) );
  EDFFX1 \rf_reg<8><31>  ( .D(n5141), .E(n5143), .CK(clk), .Q(n4854), .QN(
        n3939) );
  EDFFX1 \rf_reg<8><30>  ( .D(n5140), .E(n5143), .CK(clk), .Q(n4858), .QN(
        n3942) );
  EDFFX1 \rf_reg<8><29>  ( .D(n5139), .E(n5143), .CK(clk), .Q(n4857), .QN(
        n3949) );
  EDFFX1 \rf_reg<8><28>  ( .D(n5138), .E(n5143), .CK(clk), .Q(n4856), .QN(
        n3948) );
  EDFFX1 \rf_reg<8><27>  ( .D(n5137), .E(n5143), .CK(clk), .Q(n4855), .QN(
        n3947) );
  EDFFX1 \rf_reg<8><26>  ( .D(n5136), .E(n5143), .CK(clk), .Q(n4863), .QN(
        n3946) );
  EDFFX1 \rf_reg<8><25>  ( .D(n5135), .E(n5143), .CK(clk), .Q(n4862), .QN(
        n3945) );
  EDFFX1 \rf_reg<8><24>  ( .D(n5134), .E(n5143), .CK(clk), .Q(n4861), .QN(
        n3964) );
  EDFFX1 \rf_reg<8><23>  ( .D(n5133), .E(n5143), .CK(clk), .Q(n4860), .QN(
        n3963) );
  EDFFX1 \rf_reg<8><22>  ( .D(n5132), .E(n5143), .CK(clk), .Q(n4859), .QN(
        n3962) );
  EDFFX1 \rf_reg<8><21>  ( .D(n5131), .E(n5143), .CK(clk), .Q(n4868), .QN(
        n3961) );
  EDFFX1 \rf_reg<8><20>  ( .D(n5130), .E(n5143), .CK(clk), .Q(n4867), .QN(
        n3960) );
  EDFFX1 \rf_reg<8><19>  ( .D(n5129), .E(n5144), .CK(clk), .Q(n4866), .QN(
        n3979) );
  EDFFX1 \rf_reg<8><18>  ( .D(n5128), .E(n5144), .CK(clk), .Q(n4865), .QN(
        n3978) );
  EDFFX1 \rf_reg<8><17>  ( .D(n5127), .E(n5144), .CK(clk), .Q(n4864), .QN(
        n3977) );
  EDFFX1 \rf_reg<8><16>  ( .D(n5126), .E(n5144), .CK(clk), .Q(n4873), .QN(
        n3976) );
  EDFFX1 \rf_reg<8><15>  ( .D(n5125), .E(n5144), .CK(clk), .Q(n4872), .QN(
        n3975) );
  EDFFX1 \rf_reg<8><14>  ( .D(n5124), .E(n5144), .CK(clk), .Q(n4871), .QN(
        n3994) );
  EDFFX1 \rf_reg<8><13>  ( .D(n5123), .E(n5144), .CK(clk), .Q(n4870), .QN(
        n3993) );
  EDFFX1 \rf_reg<8><12>  ( .D(n5122), .E(n5144), .CK(clk), .Q(n4869), .QN(
        n3992) );
  EDFFX1 \rf_reg<8><11>  ( .D(n5121), .E(n5144), .CK(clk), .Q(n4879), .QN(
        n3991) );
  EDFFX1 \rf_reg<8><10>  ( .D(n5120), .E(n5144), .CK(clk), .Q(n4878), .QN(
        n3990) );
  EDFFX1 \rf_reg<8><9>  ( .D(n5119), .E(n5144), .CK(clk), .Q(n4877), .QN(n3995) );
  EDFFX1 \rf_reg<8><8>  ( .D(n5118), .E(n5144), .CK(clk), .Q(n4876), .QN(n4012) );
  EDFFX1 \rf_reg<8><7>  ( .D(n5117), .E(n1575), .CK(clk), .Q(n4875), .QN(n4011) );
  EDFFX1 \rf_reg<8><6>  ( .D(n5116), .E(n1575), .CK(clk), .Q(n4874), .QN(n4010) );
  EDFFX1 \rf_reg<8><5>  ( .D(n5115), .E(n5143), .CK(clk), .Q(n4884), .QN(n4009) );
  EDFFX1 \rf_reg<8><4>  ( .D(n5114), .E(n5144), .CK(clk), .Q(n4883), .QN(n4008) );
  EDFFX1 \rf_reg<8><3>  ( .D(n5113), .E(n5143), .CK(clk), .Q(n4882), .QN(n4026) );
  EDFFX1 \rf_reg<8><2>  ( .D(n5112), .E(n5144), .CK(clk), .Q(n4881), .QN(n4025) );
  EDFFX1 \rf_reg<8><1>  ( .D(n5111), .E(n5143), .CK(clk), .Q(n4880), .QN(n4024) );
  EDFFX1 \rf_reg<8><0>  ( .D(n5110), .E(n5144), .CK(clk), .Q(n4885), .QN(n4023) );
  EDFFX1 \rf_reg<0><31>  ( .D(n5141), .E(n5149), .CK(clk), .Q(n4981), .QN(
        n3941) );
  EDFFX1 \rf_reg<0><30>  ( .D(n5140), .E(n5149), .CK(clk), .Q(n4978), .QN(
        n3944) );
  EDFFX1 \rf_reg<0><29>  ( .D(n5139), .E(n5149), .CK(clk), .Q(n4975), .QN(
        n3959) );
  EDFFX1 \rf_reg<0><28>  ( .D(n5138), .E(n5149), .CK(clk), .Q(n4972), .QN(
        n3957) );
  EDFFX1 \rf_reg<0><27>  ( .D(n5137), .E(n5149), .CK(clk), .Q(n4969), .QN(
        n3955) );
  EDFFX1 \rf_reg<0><26>  ( .D(n5136), .E(n5149), .CK(clk), .Q(n4966), .QN(
        n3953) );
  EDFFX1 \rf_reg<0><25>  ( .D(n5135), .E(n5149), .CK(clk), .Q(n4963), .QN(
        n3951) );
  EDFFX1 \rf_reg<0><24>  ( .D(n5134), .E(n5149), .CK(clk), .Q(n4960), .QN(
        n3974) );
  EDFFX1 \rf_reg<0><23>  ( .D(n5133), .E(n5149), .CK(clk), .Q(n4957), .QN(
        n3972) );
  EDFFX1 \rf_reg<0><22>  ( .D(n5132), .E(n5149), .CK(clk), .Q(n4954), .QN(
        n3970) );
  EDFFX1 \rf_reg<0><21>  ( .D(n5131), .E(n5149), .CK(clk), .Q(n4951), .QN(
        n3968) );
  EDFFX1 \rf_reg<0><20>  ( .D(n5130), .E(n5149), .CK(clk), .Q(n4948), .QN(
        n3966) );
  EDFFX1 \rf_reg<0><19>  ( .D(n5129), .E(n5150), .CK(clk), .Q(n4945), .QN(
        n3989) );
  EDFFX1 \rf_reg<0><18>  ( .D(n5128), .E(n5150), .CK(clk), .Q(n4942), .QN(
        n3987) );
  EDFFX1 \rf_reg<0><17>  ( .D(n5127), .E(n5150), .CK(clk), .Q(n4939), .QN(
        n3985) );
  EDFFX1 \rf_reg<0><16>  ( .D(n5126), .E(n5150), .CK(clk), .Q(n4936), .QN(
        n3983) );
  EDFFX1 \rf_reg<0><15>  ( .D(n5125), .E(n5150), .CK(clk), .Q(n4933), .QN(
        n3981) );
  EDFFX1 \rf_reg<0><14>  ( .D(n5124), .E(n5150), .CK(clk), .Q(n4930), .QN(
        n4007) );
  EDFFX1 \rf_reg<0><13>  ( .D(n5123), .E(n5150), .CK(clk), .Q(n4927), .QN(
        n4005) );
  EDFFX1 \rf_reg<0><12>  ( .D(n5122), .E(n5150), .CK(clk), .Q(n4924), .QN(
        n4003) );
  EDFFX1 \rf_reg<0><11>  ( .D(n5121), .E(n5150), .CK(clk), .Q(n4921), .QN(
        n4001) );
  EDFFX1 \rf_reg<0><10>  ( .D(n5120), .E(n5150), .CK(clk), .Q(n4918), .QN(
        n3999) );
  EDFFX1 \rf_reg<0><9>  ( .D(n5119), .E(n5150), .CK(clk), .Q(n4915), .QN(n3997) );
  EDFFX1 \rf_reg<0><8>  ( .D(n5118), .E(n5150), .CK(clk), .Q(n4912), .QN(n4022) );
  EDFFX1 \rf_reg<0><7>  ( .D(n5117), .E(n1573), .CK(clk), .Q(n4909), .QN(n4020) );
  EDFFX1 \rf_reg<0><6>  ( .D(n5116), .E(n1573), .CK(clk), .Q(n4906), .QN(n4018) );
  EDFFX1 \rf_reg<0><5>  ( .D(n5115), .E(n5149), .CK(clk), .Q(n4903), .QN(n4016) );
  EDFFX1 \rf_reg<0><4>  ( .D(n5114), .E(n5150), .CK(clk), .Q(n4900), .QN(n4014) );
  EDFFX1 \rf_reg<0><3>  ( .D(n5113), .E(n5149), .CK(clk), .Q(n4897), .QN(n4034) );
  EDFFX1 \rf_reg<0><2>  ( .D(n5112), .E(n5150), .CK(clk), .Q(n4894), .QN(n4032) );
  EDFFX1 \rf_reg<0><1>  ( .D(n5111), .E(n5149), .CK(clk), .Q(n4891), .QN(n4030) );
  EDFFX1 \rf_reg<0><0>  ( .D(n5110), .E(n5150), .CK(clk), .Q(n4888), .QN(n4028) );
  EDFFX1 \rf_reg<13><31>  ( .D(n5141), .E(n5223), .CK(clk), .Q(n4755), .QN(
        n4354) );
  EDFFX1 \rf_reg<13><30>  ( .D(n5140), .E(n5223), .CK(clk), .Q(n4752), .QN(
        n4353) );
  EDFFX1 \rf_reg<13><29>  ( .D(n5139), .E(n5223), .CK(clk), .Q(n4749), .QN(
        n4352) );
  EDFFX1 \rf_reg<13><28>  ( .D(n5138), .E(n5223), .CK(clk), .Q(n4746), .QN(
        n4351) );
  EDFFX1 \rf_reg<13><27>  ( .D(n5137), .E(n5223), .CK(clk), .Q(n4743), .QN(
        n4350) );
  EDFFX1 \rf_reg<13><26>  ( .D(n5136), .E(n5223), .CK(clk), .Q(n4740), .QN(
        n4349) );
  EDFFX1 \rf_reg<13><25>  ( .D(n5135), .E(n5223), .CK(clk), .Q(n4737), .QN(
        n4348) );
  EDFFX1 \rf_reg<13><24>  ( .D(n5134), .E(n5223), .CK(clk), .Q(n4734), .QN(
        n4347) );
  EDFFX1 \rf_reg<13><23>  ( .D(n5133), .E(n5223), .CK(clk), .Q(n4731), .QN(
        n4346) );
  EDFFX1 \rf_reg<13><22>  ( .D(n5132), .E(n5223), .CK(clk), .Q(n4728), .QN(
        n4345) );
  EDFFX1 \rf_reg<13><21>  ( .D(n5131), .E(n5223), .CK(clk), .Q(n4725), .QN(
        n4344) );
  EDFFX1 \rf_reg<13><20>  ( .D(n5130), .E(n5223), .CK(clk), .Q(n4722), .QN(
        n4343) );
  EDFFX1 \rf_reg<13><19>  ( .D(n5129), .E(n5224), .CK(clk), .Q(n4719), .QN(
        n4342) );
  EDFFX1 \rf_reg<13><18>  ( .D(n5128), .E(n5224), .CK(clk), .Q(n4716), .QN(
        n4341) );
  EDFFX1 \rf_reg<13><17>  ( .D(n5127), .E(n5224), .CK(clk), .Q(n4713), .QN(
        n4340) );
  EDFFX1 \rf_reg<13><16>  ( .D(n5126), .E(n5224), .CK(clk), .Q(n4710), .QN(
        n4339) );
  EDFFX1 \rf_reg<13><15>  ( .D(n5125), .E(n5224), .CK(clk), .Q(n4707), .QN(
        n4338) );
  EDFFX1 \rf_reg<13><14>  ( .D(n5124), .E(n5224), .CK(clk), .Q(n4704), .QN(
        n4337) );
  EDFFX1 \rf_reg<13><13>  ( .D(n5123), .E(n5224), .CK(clk), .Q(n4701), .QN(
        n4336) );
  EDFFX1 \rf_reg<13><12>  ( .D(n5122), .E(n5224), .CK(clk), .Q(n4698), .QN(
        n4335) );
  EDFFX1 \rf_reg<13><11>  ( .D(n5121), .E(n5224), .CK(clk), .Q(n4695), .QN(
        n4334) );
  EDFFX1 \rf_reg<13><10>  ( .D(n5120), .E(n5224), .CK(clk), .Q(n4692), .QN(
        n4333) );
  EDFFX1 \rf_reg<13><9>  ( .D(n5119), .E(n5224), .CK(clk), .Q(n4689), .QN(
        n4332) );
  EDFFX1 \rf_reg<13><8>  ( .D(n5118), .E(n5224), .CK(clk), .Q(n4686), .QN(
        n4331) );
  EDFFX1 \rf_reg<13><7>  ( .D(n5117), .E(n5223), .CK(clk), .Q(n4683), .QN(
        n4330) );
  EDFFX1 \rf_reg<13><6>  ( .D(n5116), .E(n5224), .CK(clk), .Q(n4680), .QN(
        n4329) );
  EDFFX1 \rf_reg<13><5>  ( .D(n5115), .E(n5223), .CK(clk), .Q(n4677), .QN(
        n4328) );
  EDFFX1 \rf_reg<13><4>  ( .D(n5114), .E(n5224), .CK(clk), .Q(n4674), .QN(
        n4327) );
  EDFFX1 \rf_reg<13><3>  ( .D(n5113), .E(n5223), .CK(clk), .Q(n4671), .QN(
        n4326) );
  EDFFX1 \rf_reg<13><2>  ( .D(n5112), .E(n5224), .CK(clk), .Q(n4668), .QN(
        n4325) );
  EDFFX1 \rf_reg<13><1>  ( .D(n5111), .E(n5223), .CK(clk), .Q(n4665), .QN(
        n4324) );
  EDFFX1 \rf_reg<13><0>  ( .D(n5110), .E(n5224), .CK(clk), .Q(n4662), .QN(
        n4323) );
  EDFFX1 \rf_reg<9><31>  ( .D(n5141), .E(n5221), .CK(clk), .Q(n4630), .QN(
        n4099) );
  EDFFX1 \rf_reg<9><30>  ( .D(n5140), .E(n5221), .CK(clk), .Q(n4634), .QN(
        n4102) );
  EDFFX1 \rf_reg<9><29>  ( .D(n5139), .E(n5221), .CK(clk), .Q(n4633), .QN(
        n4109) );
  EDFFX1 \rf_reg<9><28>  ( .D(n5138), .E(n5221), .CK(clk), .Q(n4632), .QN(
        n4108) );
  EDFFX1 \rf_reg<9><27>  ( .D(n5137), .E(n5221), .CK(clk), .Q(n4631), .QN(
        n4107) );
  EDFFX1 \rf_reg<9><26>  ( .D(n5136), .E(n5221), .CK(clk), .Q(n4639), .QN(
        n4106) );
  EDFFX1 \rf_reg<9><25>  ( .D(n5135), .E(n5221), .CK(clk), .Q(n4638), .QN(
        n4105) );
  EDFFX1 \rf_reg<9><24>  ( .D(n5134), .E(n5221), .CK(clk), .Q(n4637), .QN(
        n4124) );
  EDFFX1 \rf_reg<9><23>  ( .D(n5133), .E(n5221), .CK(clk), .Q(n4636), .QN(
        n4123) );
  EDFFX1 \rf_reg<9><22>  ( .D(n5132), .E(n5221), .CK(clk), .Q(n4635), .QN(
        n4122) );
  EDFFX1 \rf_reg<9><21>  ( .D(n5131), .E(n5221), .CK(clk), .Q(n4644), .QN(
        n4121) );
  EDFFX1 \rf_reg<9><20>  ( .D(n5130), .E(n5221), .CK(clk), .Q(n4643), .QN(
        n4120) );
  EDFFX1 \rf_reg<9><19>  ( .D(n5129), .E(n5222), .CK(clk), .Q(n4642), .QN(
        n4139) );
  EDFFX1 \rf_reg<9><18>  ( .D(n5128), .E(n5222), .CK(clk), .Q(n4641), .QN(
        n4138) );
  EDFFX1 \rf_reg<9><17>  ( .D(n5127), .E(n5222), .CK(clk), .Q(n4640), .QN(
        n4137) );
  EDFFX1 \rf_reg<9><16>  ( .D(n5126), .E(n5222), .CK(clk), .Q(n4649), .QN(
        n4136) );
  EDFFX1 \rf_reg<9><15>  ( .D(n5125), .E(n5222), .CK(clk), .Q(n4648), .QN(
        n4135) );
  EDFFX1 \rf_reg<9><14>  ( .D(n5124), .E(n5222), .CK(clk), .Q(n4647), .QN(
        n4154) );
  EDFFX1 \rf_reg<9><13>  ( .D(n5123), .E(n5222), .CK(clk), .Q(n4646), .QN(
        n4153) );
  EDFFX1 \rf_reg<9><12>  ( .D(n5122), .E(n5222), .CK(clk), .Q(n4645), .QN(
        n4152) );
  EDFFX1 \rf_reg<9><11>  ( .D(n5121), .E(n5222), .CK(clk), .Q(n4655), .QN(
        n4151) );
  EDFFX1 \rf_reg<9><10>  ( .D(n5120), .E(n5222), .CK(clk), .Q(n4654), .QN(
        n4150) );
  EDFFX1 \rf_reg<9><9>  ( .D(n5119), .E(n5222), .CK(clk), .Q(n4653), .QN(n4155) );
  EDFFX1 \rf_reg<9><8>  ( .D(n5118), .E(n5222), .CK(clk), .Q(n4652), .QN(n4172) );
  EDFFX1 \rf_reg<9><7>  ( .D(n5117), .E(n5221), .CK(clk), .Q(n4651), .QN(n4171) );
  EDFFX1 \rf_reg<9><6>  ( .D(n5116), .E(n5222), .CK(clk), .Q(n4650), .QN(n4170) );
  EDFFX1 \rf_reg<9><5>  ( .D(n5115), .E(n5221), .CK(clk), .Q(n4660), .QN(n4169) );
  EDFFX1 \rf_reg<9><4>  ( .D(n5114), .E(n5222), .CK(clk), .Q(n4659), .QN(n4168) );
  EDFFX1 \rf_reg<9><3>  ( .D(n5113), .E(n5221), .CK(clk), .Q(n4658), .QN(n4186) );
  EDFFX1 \rf_reg<9><2>  ( .D(n5112), .E(n5222), .CK(clk), .Q(n4657), .QN(n4185) );
  EDFFX1 \rf_reg<9><1>  ( .D(n5111), .E(n5221), .CK(clk), .Q(n4656), .QN(n4184) );
  EDFFX1 \rf_reg<9><0>  ( .D(n5110), .E(n5222), .CK(clk), .Q(n4661), .QN(n4183) );
  EDFFX1 \rf_reg<5><31>  ( .D(n5141), .E(n5233), .CK(clk), .Q(n4756), .QN(
        n4100) );
  EDFFX1 \rf_reg<5><30>  ( .D(n5140), .E(n5233), .CK(clk), .Q(n4753), .QN(
        n4103) );
  EDFFX1 \rf_reg<5><29>  ( .D(n5139), .E(n5233), .CK(clk), .Q(n4750), .QN(
        n4118) );
  EDFFX1 \rf_reg<5><28>  ( .D(n5138), .E(n5233), .CK(clk), .Q(n4747), .QN(
        n4116) );
  EDFFX1 \rf_reg<5><27>  ( .D(n5137), .E(n5233), .CK(clk), .Q(n4744), .QN(
        n4114) );
  EDFFX1 \rf_reg<5><26>  ( .D(n5136), .E(n5233), .CK(clk), .Q(n4741), .QN(
        n4112) );
  EDFFX1 \rf_reg<5><25>  ( .D(n5135), .E(n5233), .CK(clk), .Q(n4738), .QN(
        n4110) );
  EDFFX1 \rf_reg<5><24>  ( .D(n5134), .E(n5233), .CK(clk), .Q(n4735), .QN(
        n4133) );
  EDFFX1 \rf_reg<5><23>  ( .D(n5133), .E(n5233), .CK(clk), .Q(n4732), .QN(
        n4131) );
  EDFFX1 \rf_reg<5><22>  ( .D(n5132), .E(n5233), .CK(clk), .Q(n4729), .QN(
        n4129) );
  EDFFX1 \rf_reg<5><21>  ( .D(n5131), .E(n5233), .CK(clk), .Q(n4726), .QN(
        n4127) );
  EDFFX1 \rf_reg<5><20>  ( .D(n5130), .E(n5233), .CK(clk), .Q(n4723), .QN(
        n4125) );
  EDFFX1 \rf_reg<5><19>  ( .D(n5129), .E(n5234), .CK(clk), .Q(n4720), .QN(
        n4148) );
  EDFFX1 \rf_reg<5><18>  ( .D(n5128), .E(n5234), .CK(clk), .Q(n4717), .QN(
        n4146) );
  EDFFX1 \rf_reg<5><17>  ( .D(n5127), .E(n5234), .CK(clk), .Q(n4714), .QN(
        n4144) );
  EDFFX1 \rf_reg<5><16>  ( .D(n5126), .E(n5234), .CK(clk), .Q(n4711), .QN(
        n4142) );
  EDFFX1 \rf_reg<5><15>  ( .D(n5125), .E(n5234), .CK(clk), .Q(n4708), .QN(
        n4140) );
  EDFFX1 \rf_reg<5><14>  ( .D(n5124), .E(n5234), .CK(clk), .Q(n4705), .QN(
        n4166) );
  EDFFX1 \rf_reg<5><13>  ( .D(n5123), .E(n5234), .CK(clk), .Q(n4702), .QN(
        n4164) );
  EDFFX1 \rf_reg<5><12>  ( .D(n5122), .E(n5234), .CK(clk), .Q(n4699), .QN(
        n4162) );
  EDFFX1 \rf_reg<5><11>  ( .D(n5121), .E(n5234), .CK(clk), .Q(n4696), .QN(
        n4160) );
  EDFFX1 \rf_reg<5><10>  ( .D(n5120), .E(n5234), .CK(clk), .Q(n4693), .QN(
        n4158) );
  EDFFX1 \rf_reg<5><9>  ( .D(n5119), .E(n5234), .CK(clk), .Q(n4690), .QN(n4156) );
  EDFFX1 \rf_reg<5><8>  ( .D(n5118), .E(n5234), .CK(clk), .Q(n4687), .QN(n4181) );
  EDFFX1 \rf_reg<5><7>  ( .D(n5117), .E(n5233), .CK(clk), .Q(n4684), .QN(n4179) );
  EDFFX1 \rf_reg<5><6>  ( .D(n5116), .E(n5234), .CK(clk), .Q(n4681), .QN(n4177) );
  EDFFX1 \rf_reg<5><5>  ( .D(n5115), .E(n5233), .CK(clk), .Q(n4678), .QN(n4175) );
  EDFFX1 \rf_reg<5><4>  ( .D(n5114), .E(n5234), .CK(clk), .Q(n4675), .QN(n4173) );
  EDFFX1 \rf_reg<5><3>  ( .D(n5113), .E(n5233), .CK(clk), .Q(n4672), .QN(n4193) );
  EDFFX1 \rf_reg<5><2>  ( .D(n5112), .E(n5234), .CK(clk), .Q(n4669), .QN(n4191) );
  EDFFX1 \rf_reg<5><1>  ( .D(n5111), .E(n5233), .CK(clk), .Q(n4666), .QN(n4189) );
  EDFFX1 \rf_reg<5><0>  ( .D(n5110), .E(n5234), .CK(clk), .Q(n4663), .QN(n4187) );
  EDFFX1 \rf_reg<1><31>  ( .D(n5141), .E(n5235), .CK(clk), .Q(n4757), .QN(
        n4101) );
  EDFFX1 \rf_reg<1><30>  ( .D(n5140), .E(n5235), .CK(clk), .Q(n4754), .QN(
        n4104) );
  EDFFX1 \rf_reg<1><29>  ( .D(n5139), .E(n5235), .CK(clk), .Q(n4751), .QN(
        n4119) );
  EDFFX1 \rf_reg<1><28>  ( .D(n5138), .E(n5235), .CK(clk), .Q(n4748), .QN(
        n4117) );
  EDFFX1 \rf_reg<1><27>  ( .D(n5137), .E(n5235), .CK(clk), .Q(n4745), .QN(
        n4115) );
  EDFFX1 \rf_reg<1><26>  ( .D(n5136), .E(n5235), .CK(clk), .Q(n4742), .QN(
        n4113) );
  EDFFX1 \rf_reg<1><25>  ( .D(n5135), .E(n5235), .CK(clk), .Q(n4739), .QN(
        n4111) );
  EDFFX1 \rf_reg<1><24>  ( .D(n5134), .E(n5235), .CK(clk), .Q(n4736), .QN(
        n4134) );
  EDFFX1 \rf_reg<1><23>  ( .D(n5133), .E(n5235), .CK(clk), .Q(n4733), .QN(
        n4132) );
  EDFFX1 \rf_reg<1><22>  ( .D(n5132), .E(n5235), .CK(clk), .Q(n4730), .QN(
        n4130) );
  EDFFX1 \rf_reg<1><21>  ( .D(n5131), .E(n5235), .CK(clk), .Q(n4727), .QN(
        n4128) );
  EDFFX1 \rf_reg<1><20>  ( .D(n5130), .E(n5235), .CK(clk), .Q(n4724), .QN(
        n4126) );
  EDFFX1 \rf_reg<1><19>  ( .D(n5129), .E(n5236), .CK(clk), .Q(n4721), .QN(
        n4149) );
  EDFFX1 \rf_reg<1><18>  ( .D(n5128), .E(n5236), .CK(clk), .Q(n4718), .QN(
        n4147) );
  EDFFX1 \rf_reg<1><17>  ( .D(n5127), .E(n5236), .CK(clk), .Q(n4715), .QN(
        n4145) );
  EDFFX1 \rf_reg<1><16>  ( .D(n5126), .E(n5236), .CK(clk), .Q(n4712), .QN(
        n4143) );
  EDFFX1 \rf_reg<1><15>  ( .D(n5125), .E(n5236), .CK(clk), .Q(n4709), .QN(
        n4141) );
  EDFFX1 \rf_reg<1><14>  ( .D(n5124), .E(n5236), .CK(clk), .Q(n4706), .QN(
        n4167) );
  EDFFX1 \rf_reg<1><13>  ( .D(n5123), .E(n5236), .CK(clk), .Q(n4703), .QN(
        n4165) );
  EDFFX1 \rf_reg<1><12>  ( .D(n5122), .E(n5236), .CK(clk), .Q(n4700), .QN(
        n4163) );
  EDFFX1 \rf_reg<1><11>  ( .D(n5121), .E(n5236), .CK(clk), .Q(n4697), .QN(
        n4161) );
  EDFFX1 \rf_reg<1><10>  ( .D(n5120), .E(n5236), .CK(clk), .Q(n4694), .QN(
        n4159) );
  EDFFX1 \rf_reg<1><9>  ( .D(n5119), .E(n5236), .CK(clk), .Q(n4691), .QN(n4157) );
  EDFFX1 \rf_reg<1><8>  ( .D(n5118), .E(n5236), .CK(clk), .Q(n4688), .QN(n4182) );
  EDFFX1 \rf_reg<1><7>  ( .D(n5117), .E(n5235), .CK(clk), .Q(n4685), .QN(n4180) );
  EDFFX1 \rf_reg<1><6>  ( .D(n5116), .E(n5236), .CK(clk), .Q(n4682), .QN(n4178) );
  EDFFX1 \rf_reg<1><5>  ( .D(n5115), .E(n5235), .CK(clk), .Q(n4679), .QN(n4176) );
  EDFFX1 \rf_reg<1><4>  ( .D(n5114), .E(n5236), .CK(clk), .Q(n4676), .QN(n4174) );
  EDFFX1 \rf_reg<1><3>  ( .D(n5113), .E(n5235), .CK(clk), .Q(n4673), .QN(n4194) );
  EDFFX1 \rf_reg<1><2>  ( .D(n5112), .E(n5236), .CK(clk), .Q(n4670), .QN(n4192) );
  EDFFX1 \rf_reg<1><1>  ( .D(n5111), .E(n5235), .CK(clk), .Q(n4667), .QN(n4190) );
  EDFFX1 \rf_reg<1><0>  ( .D(n5110), .E(n5236), .CK(clk), .Q(n4664), .QN(n4188) );
  EDFFX1 \rf_reg<14><31>  ( .D(n5141), .E(n5227), .CK(clk), .Q(n4386), .QN(
        n4984) );
  EDFFX1 \rf_reg<14><30>  ( .D(n5140), .E(n5227), .CK(clk), .Q(n4385), .QN(
        n4996) );
  EDFFX1 \rf_reg<14><29>  ( .D(n5139), .E(n5227), .CK(clk), .Q(n4384), .QN(
        n4993) );
  EDFFX1 \rf_reg<14><28>  ( .D(n5138), .E(n5227), .CK(clk), .Q(n4383), .QN(
        n4990) );
  EDFFX1 \rf_reg<14><27>  ( .D(n5137), .E(n5227), .CK(clk), .Q(n4382), .QN(
        n4987) );
  EDFFX1 \rf_reg<14><26>  ( .D(n5136), .E(n5227), .CK(clk), .Q(n4381), .QN(
        n5011) );
  EDFFX1 \rf_reg<14><25>  ( .D(n5135), .E(n5227), .CK(clk), .Q(n4380), .QN(
        n5008) );
  EDFFX1 \rf_reg<14><24>  ( .D(n5134), .E(n5227), .CK(clk), .Q(n4379), .QN(
        n5005) );
  EDFFX1 \rf_reg<14><23>  ( .D(n5133), .E(n5227), .CK(clk), .Q(n4378), .QN(
        n5002) );
  EDFFX1 \rf_reg<14><22>  ( .D(n5132), .E(n5227), .CK(clk), .Q(n4377), .QN(
        n4999) );
  EDFFX1 \rf_reg<14><21>  ( .D(n5131), .E(n5227), .CK(clk), .Q(n4376), .QN(
        n5026) );
  EDFFX1 \rf_reg<14><20>  ( .D(n5130), .E(n5227), .CK(clk), .Q(n4375), .QN(
        n5023) );
  EDFFX1 \rf_reg<14><19>  ( .D(n5129), .E(n5228), .CK(clk), .Q(n4374), .QN(
        n5020) );
  EDFFX1 \rf_reg<14><18>  ( .D(n5128), .E(n5228), .CK(clk), .Q(n4373), .QN(
        n5017) );
  EDFFX1 \rf_reg<14><17>  ( .D(n5127), .E(n5228), .CK(clk), .Q(n4372), .QN(
        n5014) );
  EDFFX1 \rf_reg<14><16>  ( .D(n5126), .E(n5228), .CK(clk), .Q(n4371), .QN(
        n5041) );
  EDFFX1 \rf_reg<14><15>  ( .D(n5125), .E(n5228), .CK(clk), .Q(n4370), .QN(
        n5038) );
  EDFFX1 \rf_reg<14><14>  ( .D(n5124), .E(n5228), .CK(clk), .Q(n4369), .QN(
        n5035) );
  EDFFX1 \rf_reg<14><13>  ( .D(n5123), .E(n5228), .CK(clk), .Q(n4368), .QN(
        n5032) );
  EDFFX1 \rf_reg<14><12>  ( .D(n5122), .E(n5228), .CK(clk), .Q(n4367), .QN(
        n5029) );
  EDFFX1 \rf_reg<14><11>  ( .D(n5121), .E(n5228), .CK(clk), .Q(n4366), .QN(
        n5059) );
  EDFFX1 \rf_reg<14><10>  ( .D(n5120), .E(n5228), .CK(clk), .Q(n4365), .QN(
        n5056) );
  EDFFX1 \rf_reg<14><9>  ( .D(n5119), .E(n5228), .CK(clk), .Q(n4364), .QN(
        n5053) );
  EDFFX1 \rf_reg<14><8>  ( .D(n5118), .E(n5228), .CK(clk), .Q(n4363), .QN(
        n5050) );
  EDFFX1 \rf_reg<14><7>  ( .D(n5117), .E(n1580), .CK(clk), .Q(n4362), .QN(
        n5047) );
  EDFFX1 \rf_reg<14><6>  ( .D(n5116), .E(n1580), .CK(clk), .Q(n4361), .QN(
        n5044) );
  EDFFX1 \rf_reg<14><5>  ( .D(n5115), .E(n5227), .CK(clk), .Q(n4360), .QN(
        n5074) );
  EDFFX1 \rf_reg<14><4>  ( .D(n5114), .E(n5228), .CK(clk), .Q(n4359), .QN(
        n5071) );
  EDFFX1 \rf_reg<14><3>  ( .D(n5113), .E(n5227), .CK(clk), .Q(n4358), .QN(
        n5068) );
  EDFFX1 \rf_reg<14><2>  ( .D(n5112), .E(n5228), .CK(clk), .Q(n4357), .QN(
        n5065) );
  EDFFX1 \rf_reg<14><1>  ( .D(n5111), .E(n5227), .CK(clk), .Q(n4356), .QN(
        n5062) );
  EDFFX1 \rf_reg<14><0>  ( .D(n5110), .E(n5228), .CK(clk), .Q(n4355), .QN(
        n5077) );
  EDFFX1 \rf_reg<6><31>  ( .D(n5141), .E(n5245), .CK(clk), .Q(\rf<6><31> ), 
        .QN(n4983) );
  EDFFX1 \rf_reg<6><30>  ( .D(n5140), .E(n5245), .CK(clk), .Q(\rf<6><30> ), 
        .QN(n4995) );
  EDFFX1 \rf_reg<6><29>  ( .D(n5139), .E(n5245), .CK(clk), .Q(\rf<6><29> ), 
        .QN(n4992) );
  EDFFX1 \rf_reg<6><28>  ( .D(n5138), .E(n5245), .CK(clk), .Q(\rf<6><28> ), 
        .QN(n4989) );
  EDFFX1 \rf_reg<6><27>  ( .D(n5137), .E(n5245), .CK(clk), .Q(\rf<6><27> ), 
        .QN(n4986) );
  EDFFX1 \rf_reg<6><26>  ( .D(n5136), .E(n5245), .CK(clk), .Q(\rf<6><26> ), 
        .QN(n5010) );
  EDFFX1 \rf_reg<6><25>  ( .D(n5135), .E(n5245), .CK(clk), .Q(\rf<6><25> ), 
        .QN(n5007) );
  EDFFX1 \rf_reg<6><24>  ( .D(n5134), .E(n5245), .CK(clk), .Q(\rf<6><24> ), 
        .QN(n5004) );
  EDFFX1 \rf_reg<6><23>  ( .D(n5133), .E(n5245), .CK(clk), .Q(\rf<6><23> ), 
        .QN(n5001) );
  EDFFX1 \rf_reg<6><22>  ( .D(n5132), .E(n5245), .CK(clk), .Q(\rf<6><22> ), 
        .QN(n4998) );
  EDFFX1 \rf_reg<6><21>  ( .D(n5131), .E(n5245), .CK(clk), .Q(\rf<6><21> ), 
        .QN(n5025) );
  EDFFX1 \rf_reg<6><20>  ( .D(n5130), .E(n5245), .CK(clk), .Q(\rf<6><20> ), 
        .QN(n5022) );
  EDFFX1 \rf_reg<6><19>  ( .D(n5129), .E(n5246), .CK(clk), .Q(\rf<6><19> ), 
        .QN(n5019) );
  EDFFX1 \rf_reg<6><18>  ( .D(n5128), .E(n5246), .CK(clk), .Q(\rf<6><18> ), 
        .QN(n5016) );
  EDFFX1 \rf_reg<6><17>  ( .D(n5127), .E(n5246), .CK(clk), .Q(\rf<6><17> ), 
        .QN(n5013) );
  EDFFX1 \rf_reg<6><16>  ( .D(n5126), .E(n5246), .CK(clk), .Q(\rf<6><16> ), 
        .QN(n5040) );
  EDFFX1 \rf_reg<6><15>  ( .D(n5125), .E(n5246), .CK(clk), .Q(\rf<6><15> ), 
        .QN(n5037) );
  EDFFX1 \rf_reg<6><14>  ( .D(n5124), .E(n5246), .CK(clk), .Q(\rf<6><14> ), 
        .QN(n5034) );
  EDFFX1 \rf_reg<6><13>  ( .D(n5123), .E(n5246), .CK(clk), .Q(\rf<6><13> ), 
        .QN(n5031) );
  EDFFX1 \rf_reg<6><12>  ( .D(n5122), .E(n5246), .CK(clk), .Q(\rf<6><12> ), 
        .QN(n5028) );
  EDFFX1 \rf_reg<6><11>  ( .D(n5121), .E(n5246), .CK(clk), .Q(\rf<6><11> ), 
        .QN(n5058) );
  EDFFX1 \rf_reg<6><10>  ( .D(n5120), .E(n5246), .CK(clk), .Q(\rf<6><10> ), 
        .QN(n5055) );
  EDFFX1 \rf_reg<6><9>  ( .D(n5119), .E(n5246), .CK(clk), .Q(\rf<6><9> ), .QN(
        n5052) );
  EDFFX1 \rf_reg<6><8>  ( .D(n5118), .E(n5246), .CK(clk), .Q(\rf<6><8> ), .QN(
        n5049) );
  EDFFX1 \rf_reg<6><7>  ( .D(n5117), .E(n13), .CK(clk), .Q(\rf<6><7> ), .QN(
        n5046) );
  EDFFX1 \rf_reg<6><6>  ( .D(n5116), .E(n13), .CK(clk), .Q(\rf<6><6> ), .QN(
        n5043) );
  EDFFX1 \rf_reg<6><5>  ( .D(n5115), .E(n5245), .CK(clk), .Q(\rf<6><5> ), .QN(
        n5073) );
  EDFFX1 \rf_reg<6><4>  ( .D(n5114), .E(n5246), .CK(clk), .Q(\rf<6><4> ), .QN(
        n5070) );
  EDFFX1 \rf_reg<6><3>  ( .D(n5113), .E(n5245), .CK(clk), .Q(\rf<6><3> ), .QN(
        n5067) );
  EDFFX1 \rf_reg<6><2>  ( .D(n5112), .E(n5246), .CK(clk), .Q(\rf<6><2> ), .QN(
        n5064) );
  EDFFX1 \rf_reg<6><1>  ( .D(n5111), .E(n5245), .CK(clk), .Q(\rf<6><1> ), .QN(
        n5061) );
  EDFFX1 \rf_reg<6><0>  ( .D(n5110), .E(n5246), .CK(clk), .Q(\rf<6><0> ), .QN(
        n5076) );
  EDFFX1 \rf_reg<10><31>  ( .D(n5141), .E(n5240), .CK(clk), .Q(\rf<10><31> ), 
        .QN(n5078) );
  EDFFX1 \rf_reg<10><30>  ( .D(n5140), .E(n5240), .CK(clk), .Q(\rf<10><30> ), 
        .QN(n5082) );
  EDFFX1 \rf_reg<10><29>  ( .D(n5139), .E(n5240), .CK(clk), .Q(\rf<10><29> ), 
        .QN(n5081) );
  EDFFX1 \rf_reg<10><28>  ( .D(n5138), .E(n5240), .CK(clk), .Q(\rf<10><28> ), 
        .QN(n5080) );
  EDFFX1 \rf_reg<10><27>  ( .D(n5137), .E(n5240), .CK(clk), .Q(\rf<10><27> ), 
        .QN(n5079) );
  EDFFX1 \rf_reg<10><26>  ( .D(n5136), .E(n5240), .CK(clk), .Q(\rf<10><26> ), 
        .QN(n5087) );
  EDFFX1 \rf_reg<10><25>  ( .D(n5135), .E(n5240), .CK(clk), .Q(\rf<10><25> ), 
        .QN(n5086) );
  EDFFX1 \rf_reg<10><24>  ( .D(n5134), .E(n5240), .CK(clk), .Q(\rf<10><24> ), 
        .QN(n5085) );
  EDFFX1 \rf_reg<10><23>  ( .D(n5133), .E(n5240), .CK(clk), .Q(\rf<10><23> ), 
        .QN(n5084) );
  EDFFX1 \rf_reg<10><22>  ( .D(n5132), .E(n5240), .CK(clk), .Q(\rf<10><22> ), 
        .QN(n5083) );
  EDFFX1 \rf_reg<10><21>  ( .D(n5131), .E(n5240), .CK(clk), .Q(\rf<10><21> ), 
        .QN(n5092) );
  EDFFX1 \rf_reg<10><20>  ( .D(n5130), .E(n5240), .CK(clk), .Q(\rf<10><20> ), 
        .QN(n5091) );
  EDFFX1 \rf_reg<10><19>  ( .D(n5129), .E(n5241), .CK(clk), .Q(\rf<10><19> ), 
        .QN(n5090) );
  EDFFX1 \rf_reg<10><18>  ( .D(n5128), .E(n5241), .CK(clk), .Q(\rf<10><18> ), 
        .QN(n5089) );
  EDFFX1 \rf_reg<10><17>  ( .D(n5127), .E(n5241), .CK(clk), .Q(\rf<10><17> ), 
        .QN(n5088) );
  EDFFX1 \rf_reg<10><16>  ( .D(n5126), .E(n5241), .CK(clk), .Q(\rf<10><16> ), 
        .QN(n5097) );
  EDFFX1 \rf_reg<10><15>  ( .D(n5125), .E(n5241), .CK(clk), .Q(\rf<10><15> ), 
        .QN(n5096) );
  EDFFX1 \rf_reg<10><14>  ( .D(n5124), .E(n5241), .CK(clk), .Q(\rf<10><14> ), 
        .QN(n5095) );
  EDFFX1 \rf_reg<10><13>  ( .D(n5123), .E(n5241), .CK(clk), .Q(\rf<10><13> ), 
        .QN(n5094) );
  EDFFX1 \rf_reg<10><12>  ( .D(n5122), .E(n5241), .CK(clk), .Q(\rf<10><12> ), 
        .QN(n5093) );
  EDFFX1 \rf_reg<10><11>  ( .D(n5121), .E(n5241), .CK(clk), .Q(\rf<10><11> ), 
        .QN(n5103) );
  EDFFX1 \rf_reg<10><10>  ( .D(n5120), .E(n5241), .CK(clk), .Q(\rf<10><10> ), 
        .QN(n5102) );
  EDFFX1 \rf_reg<10><9>  ( .D(n5119), .E(n5241), .CK(clk), .Q(\rf<10><9> ), 
        .QN(n5101) );
  EDFFX1 \rf_reg<10><8>  ( .D(n5118), .E(n5241), .CK(clk), .Q(\rf<10><8> ), 
        .QN(n5100) );
  EDFFX1 \rf_reg<10><7>  ( .D(n5117), .E(n15), .CK(clk), .Q(\rf<10><7> ), .QN(
        n5099) );
  EDFFX1 \rf_reg<10><6>  ( .D(n5116), .E(n15), .CK(clk), .Q(\rf<10><6> ), .QN(
        n5098) );
  EDFFX1 \rf_reg<10><5>  ( .D(n5115), .E(n5240), .CK(clk), .Q(\rf<10><5> ), 
        .QN(n5108) );
  EDFFX1 \rf_reg<10><4>  ( .D(n5114), .E(n5241), .CK(clk), .Q(\rf<10><4> ), 
        .QN(n5107) );
  EDFFX1 \rf_reg<10><3>  ( .D(n5113), .E(n5240), .CK(clk), .Q(\rf<10><3> ), 
        .QN(n5106) );
  EDFFX1 \rf_reg<10><2>  ( .D(n5112), .E(n5241), .CK(clk), .Q(\rf<10><2> ), 
        .QN(n5105) );
  EDFFX1 \rf_reg<10><1>  ( .D(n5111), .E(n5240), .CK(clk), .Q(\rf<10><1> ), 
        .QN(n5104) );
  EDFFX1 \rf_reg<10><0>  ( .D(n5110), .E(n5241), .CK(clk), .Q(\rf<10><0> ), 
        .QN(n5109) );
  EDFFX1 \rf_reg<2><31>  ( .D(n5141), .E(n5152), .CK(clk), .Q(\rf<2><31> ), 
        .QN(n4982) );
  EDFFX1 \rf_reg<2><30>  ( .D(n5140), .E(n5152), .CK(clk), .Q(\rf<2><30> ), 
        .QN(n4994) );
  EDFFX1 \rf_reg<2><29>  ( .D(n5139), .E(n5152), .CK(clk), .Q(\rf<2><29> ), 
        .QN(n4991) );
  EDFFX1 \rf_reg<2><28>  ( .D(n5138), .E(n5152), .CK(clk), .Q(\rf<2><28> ), 
        .QN(n4988) );
  EDFFX1 \rf_reg<2><27>  ( .D(n5137), .E(n5152), .CK(clk), .Q(\rf<2><27> ), 
        .QN(n4985) );
  EDFFX1 \rf_reg<2><26>  ( .D(n5136), .E(n5152), .CK(clk), .Q(\rf<2><26> ), 
        .QN(n5009) );
  EDFFX1 \rf_reg<2><25>  ( .D(n5135), .E(n5152), .CK(clk), .Q(\rf<2><25> ), 
        .QN(n5006) );
  EDFFX1 \rf_reg<2><24>  ( .D(n5134), .E(n5152), .CK(clk), .Q(\rf<2><24> ), 
        .QN(n5003) );
  EDFFX1 \rf_reg<2><23>  ( .D(n5133), .E(n5152), .CK(clk), .Q(\rf<2><23> ), 
        .QN(n5000) );
  EDFFX1 \rf_reg<2><22>  ( .D(n5132), .E(n5152), .CK(clk), .Q(\rf<2><22> ), 
        .QN(n4997) );
  EDFFX1 \rf_reg<2><21>  ( .D(n5131), .E(n5152), .CK(clk), .Q(\rf<2><21> ), 
        .QN(n5024) );
  EDFFX1 \rf_reg<2><20>  ( .D(n5130), .E(n5152), .CK(clk), .Q(\rf<2><20> ), 
        .QN(n5021) );
  EDFFX1 \rf_reg<2><19>  ( .D(n5129), .E(n5153), .CK(clk), .Q(\rf<2><19> ), 
        .QN(n5018) );
  EDFFX1 \rf_reg<2><18>  ( .D(n5128), .E(n5153), .CK(clk), .Q(\rf<2><18> ), 
        .QN(n5015) );
  EDFFX1 \rf_reg<2><17>  ( .D(n5127), .E(n5153), .CK(clk), .Q(\rf<2><17> ), 
        .QN(n5012) );
  EDFFX1 \rf_reg<2><16>  ( .D(n5126), .E(n5153), .CK(clk), .Q(\rf<2><16> ), 
        .QN(n5039) );
  EDFFX1 \rf_reg<2><15>  ( .D(n5125), .E(n5153), .CK(clk), .Q(\rf<2><15> ), 
        .QN(n5036) );
  EDFFX1 \rf_reg<2><14>  ( .D(n5124), .E(n5153), .CK(clk), .Q(\rf<2><14> ), 
        .QN(n5033) );
  EDFFX1 \rf_reg<2><13>  ( .D(n5123), .E(n5153), .CK(clk), .Q(\rf<2><13> ), 
        .QN(n5030) );
  EDFFX1 \rf_reg<2><12>  ( .D(n5122), .E(n5153), .CK(clk), .Q(\rf<2><12> ), 
        .QN(n5027) );
  EDFFX1 \rf_reg<2><11>  ( .D(n5121), .E(n5153), .CK(clk), .Q(\rf<2><11> ), 
        .QN(n5057) );
  EDFFX1 \rf_reg<2><10>  ( .D(n5120), .E(n5153), .CK(clk), .Q(\rf<2><10> ), 
        .QN(n5054) );
  EDFFX1 \rf_reg<2><9>  ( .D(n5119), .E(n5153), .CK(clk), .Q(\rf<2><9> ), .QN(
        n5051) );
  EDFFX1 \rf_reg<2><8>  ( .D(n5118), .E(n5153), .CK(clk), .Q(\rf<2><8> ), .QN(
        n5048) );
  EDFFX1 \rf_reg<2><7>  ( .D(n5117), .E(n1572), .CK(clk), .Q(\rf<2><7> ), .QN(
        n5045) );
  EDFFX1 \rf_reg<2><6>  ( .D(n5116), .E(n1572), .CK(clk), .Q(\rf<2><6> ), .QN(
        n5042) );
  EDFFX1 \rf_reg<2><5>  ( .D(n5115), .E(n5152), .CK(clk), .Q(\rf<2><5> ), .QN(
        n5072) );
  EDFFX1 \rf_reg<2><4>  ( .D(n5114), .E(n5153), .CK(clk), .Q(\rf<2><4> ), .QN(
        n5069) );
  EDFFX1 \rf_reg<2><3>  ( .D(n5113), .E(n5152), .CK(clk), .Q(\rf<2><3> ), .QN(
        n5066) );
  EDFFX1 \rf_reg<2><2>  ( .D(n5112), .E(n5153), .CK(clk), .Q(\rf<2><2> ), .QN(
        n5063) );
  EDFFX1 \rf_reg<2><1>  ( .D(n5111), .E(n5152), .CK(clk), .Q(\rf<2><1> ), .QN(
        n5060) );
  EDFFX1 \rf_reg<2><0>  ( .D(n5110), .E(n5153), .CK(clk), .Q(\rf<2><0> ), .QN(
        n5075) );
  EDFFX1 \rf_reg<3><31>  ( .D(n5141), .E(n5225), .CK(clk), .Q(n4418), .QN(
        n4760) );
  EDFFX1 \rf_reg<3><30>  ( .D(n5140), .E(n5225), .CK(clk), .Q(n4417), .QN(
        n4772) );
  EDFFX1 \rf_reg<3><29>  ( .D(n5139), .E(n5225), .CK(clk), .Q(n4416), .QN(
        n4769) );
  EDFFX1 \rf_reg<3><28>  ( .D(n5138), .E(n5225), .CK(clk), .Q(n4415), .QN(
        n4766) );
  EDFFX1 \rf_reg<3><27>  ( .D(n5137), .E(n5225), .CK(clk), .Q(n4414), .QN(
        n4763) );
  EDFFX1 \rf_reg<3><26>  ( .D(n5136), .E(n5225), .CK(clk), .Q(n4413), .QN(
        n4787) );
  EDFFX1 \rf_reg<3><25>  ( .D(n5135), .E(n5225), .CK(clk), .Q(n4412), .QN(
        n4784) );
  EDFFX1 \rf_reg<3><24>  ( .D(n5134), .E(n5225), .CK(clk), .Q(n4411), .QN(
        n4781) );
  EDFFX1 \rf_reg<3><23>  ( .D(n5133), .E(n5225), .CK(clk), .Q(n4410), .QN(
        n4778) );
  EDFFX1 \rf_reg<3><22>  ( .D(n5132), .E(n5225), .CK(clk), .Q(n4409), .QN(
        n4775) );
  EDFFX1 \rf_reg<3><21>  ( .D(n5131), .E(n5225), .CK(clk), .Q(n4408), .QN(
        n4802) );
  EDFFX1 \rf_reg<3><20>  ( .D(n5130), .E(n5225), .CK(clk), .Q(n4407), .QN(
        n4799) );
  EDFFX1 \rf_reg<3><19>  ( .D(n5129), .E(n5226), .CK(clk), .Q(n4406), .QN(
        n4796) );
  EDFFX1 \rf_reg<3><18>  ( .D(n5128), .E(n5226), .CK(clk), .Q(n4405), .QN(
        n4793) );
  EDFFX1 \rf_reg<3><17>  ( .D(n5127), .E(n5226), .CK(clk), .Q(n4404), .QN(
        n4790) );
  EDFFX1 \rf_reg<3><16>  ( .D(n5126), .E(n5226), .CK(clk), .Q(n4403), .QN(
        n4817) );
  EDFFX1 \rf_reg<3><15>  ( .D(n5125), .E(n5226), .CK(clk), .Q(n4402), .QN(
        n4814) );
  EDFFX1 \rf_reg<3><14>  ( .D(n5124), .E(n5226), .CK(clk), .Q(n4401), .QN(
        n4811) );
  EDFFX1 \rf_reg<3><13>  ( .D(n5123), .E(n5226), .CK(clk), .Q(n4400), .QN(
        n4808) );
  EDFFX1 \rf_reg<3><12>  ( .D(n5122), .E(n5226), .CK(clk), .Q(n4399), .QN(
        n4805) );
  EDFFX1 \rf_reg<3><11>  ( .D(n5121), .E(n5226), .CK(clk), .Q(n4398), .QN(
        n4835) );
  EDFFX1 \rf_reg<3><10>  ( .D(n5120), .E(n5226), .CK(clk), .Q(n4397), .QN(
        n4832) );
  EDFFX1 \rf_reg<3><9>  ( .D(n5119), .E(n5226), .CK(clk), .Q(n4396), .QN(n4829) );
  EDFFX1 \rf_reg<3><8>  ( .D(n5118), .E(n5226), .CK(clk), .Q(n4395), .QN(n4826) );
  EDFFX1 \rf_reg<3><7>  ( .D(n5117), .E(n5225), .CK(clk), .Q(n4394), .QN(n4823) );
  EDFFX1 \rf_reg<3><6>  ( .D(n5116), .E(n5226), .CK(clk), .Q(n4393), .QN(n4820) );
  EDFFX1 \rf_reg<3><5>  ( .D(n5115), .E(n5225), .CK(clk), .Q(n4392), .QN(n4850) );
  EDFFX1 \rf_reg<3><4>  ( .D(n5114), .E(n5226), .CK(clk), .Q(n4391), .QN(n4847) );
  EDFFX1 \rf_reg<3><3>  ( .D(n5113), .E(n5225), .CK(clk), .Q(n4390), .QN(n4844) );
  EDFFX1 \rf_reg<3><2>  ( .D(n5112), .E(n5226), .CK(clk), .Q(n4389), .QN(n4841) );
  EDFFX1 \rf_reg<3><1>  ( .D(n5111), .E(n5225), .CK(clk), .Q(n4388), .QN(n4838) );
  EDFFX1 \rf_reg<3><0>  ( .D(n5110), .E(n5226), .CK(clk), .Q(n4387), .QN(n4853) );
  EDFFX1 \rf_reg<11><31>  ( .D(n5141), .E(n16), .CK(clk), .Q(\rf<11><31> ), 
        .QN(n4759) );
  EDFFX1 \rf_reg<11><30>  ( .D(n5140), .E(n5237), .CK(clk), .Q(\rf<11><30> ), 
        .QN(n4771) );
  EDFFX1 \rf_reg<11><29>  ( .D(n5139), .E(n5238), .CK(clk), .Q(\rf<11><29> ), 
        .QN(n4768) );
  EDFFX1 \rf_reg<11><28>  ( .D(n5138), .E(n5237), .CK(clk), .Q(\rf<11><28> ), 
        .QN(n4765) );
  EDFFX1 \rf_reg<11><27>  ( .D(n5137), .E(n5238), .CK(clk), .Q(\rf<11><27> ), 
        .QN(n4762) );
  EDFFX1 \rf_reg<11><26>  ( .D(n5136), .E(n5237), .CK(clk), .Q(\rf<11><26> ), 
        .QN(n4786) );
  EDFFX1 \rf_reg<11><25>  ( .D(n5135), .E(n5238), .CK(clk), .Q(\rf<11><25> ), 
        .QN(n4783) );
  EDFFX1 \rf_reg<11><24>  ( .D(n5134), .E(n5237), .CK(clk), .Q(\rf<11><24> ), 
        .QN(n4780) );
  EDFFX1 \rf_reg<11><23>  ( .D(n5133), .E(n5238), .CK(clk), .Q(\rf<11><23> ), 
        .QN(n4777) );
  EDFFX1 \rf_reg<11><22>  ( .D(n5132), .E(n5238), .CK(clk), .Q(\rf<11><22> ), 
        .QN(n4774) );
  EDFFX1 \rf_reg<11><21>  ( .D(n5131), .E(n5238), .CK(clk), .Q(\rf<11><21> ), 
        .QN(n4801) );
  EDFFX1 \rf_reg<11><20>  ( .D(n5130), .E(n5238), .CK(clk), .Q(\rf<11><20> ), 
        .QN(n4798) );
  EDFFX1 \rf_reg<11><19>  ( .D(n5129), .E(n5237), .CK(clk), .Q(\rf<11><19> ), 
        .QN(n4795) );
  EDFFX1 \rf_reg<11><18>  ( .D(n5128), .E(n5237), .CK(clk), .Q(\rf<11><18> ), 
        .QN(n4792) );
  EDFFX1 \rf_reg<11><17>  ( .D(n5127), .E(n5237), .CK(clk), .Q(\rf<11><17> ), 
        .QN(n4789) );
  EDFFX1 \rf_reg<11><16>  ( .D(n5126), .E(n5237), .CK(clk), .Q(\rf<11><16> ), 
        .QN(n4816) );
  EDFFX1 \rf_reg<11><15>  ( .D(n5125), .E(n5237), .CK(clk), .Q(\rf<11><15> ), 
        .QN(n4813) );
  EDFFX1 \rf_reg<11><14>  ( .D(n5124), .E(n5237), .CK(clk), .Q(\rf<11><14> ), 
        .QN(n4810) );
  EDFFX1 \rf_reg<11><13>  ( .D(n5123), .E(n5237), .CK(clk), .Q(\rf<11><13> ), 
        .QN(n4807) );
  EDFFX1 \rf_reg<11><12>  ( .D(n5122), .E(n5237), .CK(clk), .Q(\rf<11><12> ), 
        .QN(n4804) );
  EDFFX1 \rf_reg<11><11>  ( .D(n5121), .E(n5237), .CK(clk), .Q(\rf<11><11> ), 
        .QN(n4834) );
  EDFFX1 \rf_reg<11><10>  ( .D(n5120), .E(n5237), .CK(clk), .Q(\rf<11><10> ), 
        .QN(n4831) );
  EDFFX1 \rf_reg<11><9>  ( .D(n5119), .E(n5237), .CK(clk), .Q(\rf<11><9> ), 
        .QN(n4828) );
  EDFFX1 \rf_reg<11><8>  ( .D(n5118), .E(n5237), .CK(clk), .Q(\rf<11><8> ), 
        .QN(n4825) );
  EDFFX1 \rf_reg<11><7>  ( .D(n5117), .E(n5238), .CK(clk), .Q(\rf<11><7> ), 
        .QN(n4822) );
  EDFFX1 \rf_reg<11><6>  ( .D(n5116), .E(n5238), .CK(clk), .Q(\rf<11><6> ), 
        .QN(n4819) );
  EDFFX1 \rf_reg<11><5>  ( .D(n5115), .E(n5238), .CK(clk), .Q(\rf<11><5> ), 
        .QN(n4849) );
  EDFFX1 \rf_reg<11><4>  ( .D(n5114), .E(n5238), .CK(clk), .Q(\rf<11><4> ), 
        .QN(n4846) );
  EDFFX1 \rf_reg<11><3>  ( .D(n5113), .E(n5238), .CK(clk), .Q(\rf<11><3> ), 
        .QN(n4843) );
  EDFFX1 \rf_reg<11><2>  ( .D(n5112), .E(n5238), .CK(clk), .Q(\rf<11><2> ), 
        .QN(n4840) );
  EDFFX1 \rf_reg<11><1>  ( .D(n5111), .E(n5238), .CK(clk), .Q(\rf<11><1> ), 
        .QN(n4837) );
  EDFFX1 \rf_reg<11><0>  ( .D(n5110), .E(n5238), .CK(clk), .Q(\rf<11><0> ), 
        .QN(n4852) );
  EDFFX1 \rf_reg<7><31>  ( .D(n5141), .E(n5243), .CK(clk), .Q(\rf<7><31> ), 
        .QN(n4758) );
  EDFFX1 \rf_reg<7><30>  ( .D(n5140), .E(n5243), .CK(clk), .Q(\rf<7><30> ), 
        .QN(n4770) );
  EDFFX1 \rf_reg<7><29>  ( .D(n5139), .E(n5243), .CK(clk), .Q(\rf<7><29> ), 
        .QN(n4767) );
  EDFFX1 \rf_reg<7><28>  ( .D(n5138), .E(n5243), .CK(clk), .Q(\rf<7><28> ), 
        .QN(n4764) );
  EDFFX1 \rf_reg<7><27>  ( .D(n5137), .E(n5243), .CK(clk), .Q(\rf<7><27> ), 
        .QN(n4761) );
  EDFFX1 \rf_reg<7><26>  ( .D(n5136), .E(n5243), .CK(clk), .Q(\rf<7><26> ), 
        .QN(n4785) );
  EDFFX1 \rf_reg<7><25>  ( .D(n5135), .E(n5243), .CK(clk), .Q(\rf<7><25> ), 
        .QN(n4782) );
  EDFFX1 \rf_reg<7><24>  ( .D(n5134), .E(n5243), .CK(clk), .Q(\rf<7><24> ), 
        .QN(n4779) );
  EDFFX1 \rf_reg<7><23>  ( .D(n5133), .E(n5243), .CK(clk), .Q(\rf<7><23> ), 
        .QN(n4776) );
  EDFFX1 \rf_reg<7><22>  ( .D(n5132), .E(n5243), .CK(clk), .Q(\rf<7><22> ), 
        .QN(n4773) );
  EDFFX1 \rf_reg<7><21>  ( .D(n5131), .E(n5243), .CK(clk), .Q(\rf<7><21> ), 
        .QN(n4800) );
  EDFFX1 \rf_reg<7><20>  ( .D(n5130), .E(n5243), .CK(clk), .Q(\rf<7><20> ), 
        .QN(n4797) );
  EDFFX1 \rf_reg<7><19>  ( .D(n5129), .E(n5244), .CK(clk), .Q(\rf<7><19> ), 
        .QN(n4794) );
  EDFFX1 \rf_reg<7><18>  ( .D(n5128), .E(n5244), .CK(clk), .Q(\rf<7><18> ), 
        .QN(n4791) );
  EDFFX1 \rf_reg<7><17>  ( .D(n5127), .E(n5244), .CK(clk), .Q(\rf<7><17> ), 
        .QN(n4788) );
  EDFFX1 \rf_reg<7><16>  ( .D(n5126), .E(n5244), .CK(clk), .Q(\rf<7><16> ), 
        .QN(n4815) );
  EDFFX1 \rf_reg<7><15>  ( .D(n5125), .E(n5244), .CK(clk), .Q(\rf<7><15> ), 
        .QN(n4812) );
  EDFFX1 \rf_reg<7><14>  ( .D(n5124), .E(n5244), .CK(clk), .Q(\rf<7><14> ), 
        .QN(n4809) );
  EDFFX1 \rf_reg<7><13>  ( .D(n5123), .E(n5244), .CK(clk), .Q(\rf<7><13> ), 
        .QN(n4806) );
  EDFFX1 \rf_reg<7><12>  ( .D(n5122), .E(n5244), .CK(clk), .Q(\rf<7><12> ), 
        .QN(n4803) );
  EDFFX1 \rf_reg<7><11>  ( .D(n5121), .E(n5244), .CK(clk), .Q(\rf<7><11> ), 
        .QN(n4833) );
  EDFFX1 \rf_reg<7><10>  ( .D(n5120), .E(n5244), .CK(clk), .Q(\rf<7><10> ), 
        .QN(n4830) );
  EDFFX1 \rf_reg<7><9>  ( .D(n5119), .E(n5244), .CK(clk), .Q(\rf<7><9> ), .QN(
        n4827) );
  EDFFX1 \rf_reg<7><8>  ( .D(n5118), .E(n5244), .CK(clk), .Q(\rf<7><8> ), .QN(
        n4824) );
  EDFFX1 \rf_reg<7><7>  ( .D(n5117), .E(n5243), .CK(clk), .Q(\rf<7><7> ), .QN(
        n4821) );
  EDFFX1 \rf_reg<7><6>  ( .D(n5116), .E(n5244), .CK(clk), .Q(\rf<7><6> ), .QN(
        n4818) );
  EDFFX1 \rf_reg<7><5>  ( .D(n5115), .E(n5243), .CK(clk), .Q(\rf<7><5> ), .QN(
        n4848) );
  EDFFX1 \rf_reg<7><4>  ( .D(n5114), .E(n5244), .CK(clk), .Q(\rf<7><4> ), .QN(
        n4845) );
  EDFFX1 \rf_reg<7><3>  ( .D(n5113), .E(n5243), .CK(clk), .Q(\rf<7><3> ), .QN(
        n4842) );
  EDFFX1 \rf_reg<7><2>  ( .D(n5112), .E(n5244), .CK(clk), .Q(\rf<7><2> ), .QN(
        n4839) );
  EDFFX1 \rf_reg<7><1>  ( .D(n5111), .E(n5243), .CK(clk), .Q(\rf<7><1> ), .QN(
        n4836) );
  EDFFX1 \rf_reg<7><0>  ( .D(n5110), .E(n5244), .CK(clk), .Q(\rf<7><0> ), .QN(
        n4851) );
  AND2X2 U4 ( .A(n1278), .B(n5288), .Y(n4602) );
  NAND2X1 U5 ( .A(n1277), .B(n5142), .Y(n4603) );
  NAND3X1 U6 ( .A(n5142), .B(n5290), .C(n1281), .Y(n4604) );
  NAND2X1 U7 ( .A(n1277), .B(n5288), .Y(n4605) );
  NAND3X1 U8 ( .A(n5288), .B(n5290), .C(n1281), .Y(n4606) );
  AND3X2 U9 ( .A(n1281), .B(n5142), .C(N17), .Y(n4607) );
  AND3X2 U10 ( .A(n1279), .B(n5142), .C(N19), .Y(n4608) );
  AND3X2 U11 ( .A(n1281), .B(n5288), .C(N17), .Y(n4609) );
  AND3X2 U12 ( .A(n5142), .B(n5286), .C(n1279), .Y(n4610) );
  AND3X2 U13 ( .A(n5288), .B(n5286), .C(n1279), .Y(n4611) );
  AND2X2 U14 ( .A(n1278), .B(n5142), .Y(n4612) );
  NAND4XL U15 ( .A(n5142), .B(n5290), .C(n5284), .D(n5286), .Y(n4613) );
  NAND4X1 U16 ( .A(n5288), .B(n5290), .C(n5284), .D(n5286), .Y(n4614) );
  AND2X2 U17 ( .A(n1562), .B(n1558), .Y(n4615) );
  AND2X2 U18 ( .A(n1558), .B(n1560), .Y(n4616) );
  AND2X2 U19 ( .A(n1558), .B(n1555), .Y(n4617) );
  AND2X2 U20 ( .A(n1553), .B(n1558), .Y(n4618) );
  AND2X2 U21 ( .A(n1557), .B(n1560), .Y(n4619) );
  AND2X2 U22 ( .A(n1557), .B(n1555), .Y(n4620) );
  AND2X2 U23 ( .A(n1553), .B(n1557), .Y(n4621) );
  OR2X2 U24 ( .A(n1566), .B(n1569), .Y(n4622) );
  OR2X2 U25 ( .A(n1567), .B(n1569), .Y(n4623) );
  NAND4X1 U26 ( .A(N19), .B(n5142), .C(n5290), .D(n5284), .Y(n4624) );
  OR2X2 U27 ( .A(n1570), .B(n1571), .Y(n4625) );
  OR2X2 U28 ( .A(n1565), .B(n1570), .Y(n4626) );
  NAND4X1 U29 ( .A(N19), .B(n5288), .C(n5290), .D(n5284), .Y(n4627) );
  OR2X2 U30 ( .A(n1566), .B(n1570), .Y(n4628) );
  OR2X2 U31 ( .A(n1567), .B(n1570), .Y(n4629) );
  INVX1 U32 ( .A(N18), .Y(n5284) );
  CLKINVX3 U33 ( .A(n5158), .Y(n5157) );
  CLKINVX3 U34 ( .A(n5183), .Y(n5182) );
  CLKINVX3 U35 ( .A(n5167), .Y(n5166) );
  CLKINVX3 U36 ( .A(n4605), .Y(n5214) );
  CLKINVX3 U37 ( .A(n4606), .Y(n5198) );
  CLKINVX3 U38 ( .A(n4614), .Y(n5206) );
  CLKINVX3 U39 ( .A(n5156), .Y(n5155) );
  CLKINVX3 U40 ( .A(n5173), .Y(n5172) );
  CLKINVX3 U41 ( .A(n4615), .Y(n5163) );
  CLKINVX3 U42 ( .A(n4618), .Y(n5187) );
  CLKINVX3 U43 ( .A(n4617), .Y(n5179) );
  CLKINVX3 U44 ( .A(n4616), .Y(n5171) );
  CLKINVX3 U45 ( .A(n5161), .Y(n5159) );
  CLKINVX3 U46 ( .A(n4621), .Y(n5185) );
  CLKINVX3 U47 ( .A(n4620), .Y(n5177) );
  CLKINVX3 U48 ( .A(n4619), .Y(n5169) );
  CLKINVX3 U49 ( .A(n4602), .Y(n5218) );
  CLKINVX3 U50 ( .A(n4611), .Y(n5210) );
  CLKINVX3 U51 ( .A(n5151), .Y(n5150) );
  INVX1 U52 ( .A(n5161), .Y(n5160) );
  CLKINVX3 U53 ( .A(n4624), .Y(n5190) );
  INVX1 U54 ( .A(n1291), .Y(n5183) );
  CLKINVX3 U55 ( .A(n5175), .Y(n5174) );
  INVX1 U56 ( .A(n1296), .Y(n5175) );
  CLKINVX3 U57 ( .A(n4627), .Y(n5189) );
  CLKINVX3 U58 ( .A(n4605), .Y(n5213) );
  CLKINVX3 U59 ( .A(n4606), .Y(n5197) );
  CLKINVX3 U60 ( .A(n4614), .Y(n5205) );
  INVX1 U61 ( .A(n1307), .Y(n5156) );
  CLKINVX3 U62 ( .A(n5181), .Y(n5180) );
  INVX1 U63 ( .A(n1292), .Y(n5181) );
  INVX1 U64 ( .A(n1297), .Y(n5173) );
  CLKINVX3 U65 ( .A(n5165), .Y(n5164) );
  INVX1 U66 ( .A(n1302), .Y(n5165) );
  CLKINVX3 U67 ( .A(n4617), .Y(n5178) );
  CLKINVX3 U68 ( .A(n4616), .Y(n5170) );
  CLKINVX3 U69 ( .A(n4621), .Y(n5184) );
  CLKINVX3 U70 ( .A(n4620), .Y(n5176) );
  CLKINVX3 U71 ( .A(n4619), .Y(n5168) );
  CLKINVX3 U72 ( .A(n4612), .Y(n5196) );
  CLKINVX3 U73 ( .A(n4610), .Y(n5219) );
  CLKINVX3 U74 ( .A(n4608), .Y(n5203) );
  CLKINVX3 U75 ( .A(n4607), .Y(n5211) );
  CLKINVX3 U76 ( .A(n5194), .Y(n5193) );
  CLKINVX3 U77 ( .A(n4609), .Y(n5202) );
  CLKINVX3 U78 ( .A(n4611), .Y(n5209) );
  CLKINVX3 U79 ( .A(n5154), .Y(n5153) );
  CLKINVX3 U80 ( .A(n5242), .Y(n5241) );
  CLKINVX3 U81 ( .A(n5145), .Y(n5144) );
  CLKINVX3 U82 ( .A(n4625), .Y(n5244) );
  CLKINVX3 U83 ( .A(n5239), .Y(n5237) );
  CLKINVX3 U84 ( .A(n4628), .Y(n5236) );
  CLKINVX3 U85 ( .A(n4629), .Y(n5234) );
  CLKINVX3 U86 ( .A(n4622), .Y(n5222) );
  CLKINVX3 U87 ( .A(n5232), .Y(n5231) );
  CLKINVX3 U88 ( .A(n4623), .Y(n5224) );
  CLKINVX3 U89 ( .A(n5247), .Y(n5246) );
  CLKINVX3 U90 ( .A(n5148), .Y(n5147) );
  CLKINVX3 U91 ( .A(n5229), .Y(n5228) );
  CLKINVX3 U92 ( .A(n4626), .Y(n5226) );
  CLKINVX3 U93 ( .A(n5151), .Y(n5149) );
  INVX1 U94 ( .A(n1573), .Y(n5151) );
  CLKINVX3 U95 ( .A(n4624), .Y(n5191) );
  CLKINVX3 U96 ( .A(n4603), .Y(n5216) );
  CLKINVX3 U97 ( .A(n4604), .Y(n5200) );
  CLKINVX3 U98 ( .A(n4613), .Y(n5208) );
  CLKINVX3 U99 ( .A(n4610), .Y(n5220) );
  CLKINVX3 U100 ( .A(n4608), .Y(n5204) );
  CLKINVX3 U101 ( .A(n4607), .Y(n5212) );
  CLKINVX3 U102 ( .A(n5239), .Y(n5238) );
  INVX1 U103 ( .A(n1304), .Y(n5161) );
  INVX1 U104 ( .A(n1306), .Y(n5158) );
  INVX1 U105 ( .A(n1301), .Y(n5167) );
  CLKINVX3 U106 ( .A(n4615), .Y(n5162) );
  CLKINVX3 U107 ( .A(n4618), .Y(n5186) );
  CLKINVX3 U108 ( .A(n4602), .Y(n5217) );
  NOR2X1 U109 ( .A(n5280), .B(n5281), .Y(n1553) );
  NOR3X1 U110 ( .A(n5290), .B(n5284), .C(n5286), .Y(n1278) );
  NOR2X1 U111 ( .A(n1564), .B(n1566), .Y(n1573) );
  NAND2X1 U112 ( .A(n1562), .B(n1557), .Y(n1304) );
  AND2X2 U113 ( .A(n1554), .B(n1560), .Y(n1302) );
  AND2X2 U114 ( .A(n1562), .B(n1554), .Y(n1307) );
  AND2X2 U115 ( .A(n1553), .B(n1556), .Y(n1306) );
  AND2X2 U116 ( .A(n1553), .B(n1554), .Y(n1292) );
  AND2X2 U117 ( .A(n1562), .B(n1556), .Y(n1301) );
  AND2X2 U118 ( .A(n1560), .B(n1556), .Y(n1296) );
  AND2X2 U119 ( .A(n1555), .B(n1556), .Y(n1291) );
  AND2X2 U120 ( .A(n1555), .B(n1554), .Y(n1297) );
  CLKINVX3 U121 ( .A(n4603), .Y(n5215) );
  CLKINVX3 U122 ( .A(n4604), .Y(n5199) );
  CLKINVX3 U123 ( .A(n4613), .Y(n5207) );
  CLKINVX3 U124 ( .A(n4627), .Y(n5188) );
  CLKINVX3 U125 ( .A(n5194), .Y(n5192) );
  INVX1 U126 ( .A(n1028), .Y(n5194) );
  CLKINVX3 U127 ( .A(n4609), .Y(n5201) );
  CLKINVX3 U128 ( .A(n5154), .Y(n5152) );
  INVX1 U129 ( .A(n1572), .Y(n5154) );
  CLKINVX3 U130 ( .A(n5242), .Y(n5240) );
  INVX1 U131 ( .A(n15), .Y(n5242) );
  CLKINVX3 U132 ( .A(n5145), .Y(n5143) );
  INVX1 U133 ( .A(n1575), .Y(n5145) );
  CLKINVX3 U134 ( .A(n4625), .Y(n5243) );
  CLKINVX3 U135 ( .A(n4628), .Y(n5235) );
  CLKINVX3 U136 ( .A(n4629), .Y(n5233) );
  CLKINVX3 U137 ( .A(n4622), .Y(n5221) );
  CLKINVX3 U138 ( .A(n5232), .Y(n5230) );
  INVX1 U139 ( .A(n1579), .Y(n5232) );
  CLKINVX3 U140 ( .A(n4623), .Y(n5223) );
  CLKINVX3 U141 ( .A(n5247), .Y(n5245) );
  INVX1 U142 ( .A(n13), .Y(n5247) );
  CLKINVX3 U143 ( .A(n5148), .Y(n5146) );
  INVX1 U144 ( .A(n1574), .Y(n5148) );
  CLKINVX3 U145 ( .A(n5229), .Y(n5227) );
  INVX1 U146 ( .A(n1580), .Y(n5229) );
  CLKINVX3 U147 ( .A(n4626), .Y(n5225) );
  INVX1 U148 ( .A(n16), .Y(n5239) );
  CLKINVX3 U149 ( .A(n4612), .Y(n5195) );
  BUFX3 U150 ( .A(\wd3<31> ), .Y(n5141) );
  OR4X2 U151 ( .A(n1080), .B(n1081), .C(n1082), .D(n1083), .Y(\rd2<31> ) );
  OAI221XL U152 ( .A0(n5212), .A1(n4758), .B0(n5210), .B1(n4982), .C0(n1085), 
        .Y(n1082) );
  OAI221XL U153 ( .A0(n5204), .A1(n4759), .B0(n5202), .B1(n4983), .C0(n1086), 
        .Y(n1081) );
  OAI221XL U154 ( .A0(n5220), .A1(n4760), .B0(n5218), .B1(n4984), .C0(n1084), 
        .Y(n1083) );
  BUFX3 U155 ( .A(\wd3<28> ), .Y(n5138) );
  BUFX3 U156 ( .A(\wd3<29> ), .Y(n5139) );
  BUFX3 U157 ( .A(\wd3<30> ), .Y(n5140) );
  OR4X2 U158 ( .A(n1120), .B(n1121), .C(n1122), .D(n1123), .Y(\rd2<27> ) );
  OAI221XL U159 ( .A0(n5211), .A1(n4761), .B0(n5210), .B1(n4985), .C0(n1125), 
        .Y(n1122) );
  OAI221XL U160 ( .A0(n5203), .A1(n4762), .B0(n5202), .B1(n4986), .C0(n1126), 
        .Y(n1121) );
  OAI221XL U161 ( .A0(n5219), .A1(n4763), .B0(n5218), .B1(n4987), .C0(n1124), 
        .Y(n1123) );
  OR4X2 U162 ( .A(n1112), .B(n1113), .C(n1114), .D(n1115), .Y(\rd2<28> ) );
  OAI221XL U163 ( .A0(n5211), .A1(n4764), .B0(n5210), .B1(n4988), .C0(n1117), 
        .Y(n1114) );
  OAI221XL U164 ( .A0(n5203), .A1(n4765), .B0(n5202), .B1(n4989), .C0(n1118), 
        .Y(n1113) );
  OAI221XL U165 ( .A0(n5219), .A1(n4766), .B0(n5218), .B1(n4990), .C0(n1116), 
        .Y(n1115) );
  OR4X2 U166 ( .A(n1104), .B(n1105), .C(n1106), .D(n1107), .Y(\rd2<29> ) );
  OAI221XL U167 ( .A0(n5211), .A1(n4767), .B0(n5210), .B1(n4991), .C0(n1109), 
        .Y(n1106) );
  OAI221XL U168 ( .A0(n5203), .A1(n4768), .B0(n5202), .B1(n4992), .C0(n1110), 
        .Y(n1105) );
  OAI221XL U169 ( .A0(n5219), .A1(n4769), .B0(n5218), .B1(n4993), .C0(n1108), 
        .Y(n1107) );
  OR4X2 U170 ( .A(n1088), .B(n1089), .C(n1090), .D(n1091), .Y(\rd2<30> ) );
  OAI221XL U171 ( .A0(n5211), .A1(n4770), .B0(n5210), .B1(n4994), .C0(n1093), 
        .Y(n1090) );
  OAI221XL U172 ( .A0(n5203), .A1(n4771), .B0(n5202), .B1(n4995), .C0(n1094), 
        .Y(n1089) );
  OAI221XL U173 ( .A0(n5219), .A1(n4772), .B0(n5218), .B1(n4996), .C0(n1092), 
        .Y(n1091) );
  BUFX3 U174 ( .A(\wd3<23> ), .Y(n5133) );
  BUFX3 U175 ( .A(\wd3<24> ), .Y(n5134) );
  BUFX3 U176 ( .A(\wd3<25> ), .Y(n5135) );
  BUFX3 U177 ( .A(\wd3<26> ), .Y(n5136) );
  BUFX3 U178 ( .A(\wd3<27> ), .Y(n5137) );
  OR4X2 U179 ( .A(n1160), .B(n1161), .C(n1162), .D(n1163), .Y(\rd2<22> ) );
  OAI221XL U180 ( .A0(n5211), .A1(n4773), .B0(n5210), .B1(n4997), .C0(n1165), 
        .Y(n1162) );
  OAI221XL U181 ( .A0(n5203), .A1(n4774), .B0(n5202), .B1(n4998), .C0(n1166), 
        .Y(n1161) );
  OAI221XL U182 ( .A0(n5219), .A1(n4775), .B0(n5218), .B1(n4999), .C0(n1164), 
        .Y(n1163) );
  OR4X2 U183 ( .A(n1152), .B(n1153), .C(n1154), .D(n1155), .Y(\rd2<23> ) );
  OAI221XL U184 ( .A0(n5211), .A1(n4776), .B0(n5210), .B1(n5000), .C0(n1157), 
        .Y(n1154) );
  OAI221XL U185 ( .A0(n5203), .A1(n4777), .B0(n5202), .B1(n5001), .C0(n1158), 
        .Y(n1153) );
  OAI221XL U186 ( .A0(n5219), .A1(n4778), .B0(n5218), .B1(n5002), .C0(n1156), 
        .Y(n1155) );
  OR4X2 U187 ( .A(n1144), .B(n1145), .C(n1146), .D(n1147), .Y(\rd2<24> ) );
  OAI221XL U188 ( .A0(n5211), .A1(n4779), .B0(n5210), .B1(n5003), .C0(n1149), 
        .Y(n1146) );
  OAI221XL U189 ( .A0(n5203), .A1(n4780), .B0(n5202), .B1(n5004), .C0(n1150), 
        .Y(n1145) );
  OAI221XL U190 ( .A0(n5219), .A1(n4781), .B0(n5218), .B1(n5005), .C0(n1148), 
        .Y(n1147) );
  OR4X2 U191 ( .A(n1136), .B(n1137), .C(n1138), .D(n1139), .Y(\rd2<25> ) );
  OAI221XL U192 ( .A0(n5211), .A1(n4782), .B0(n5210), .B1(n5006), .C0(n1141), 
        .Y(n1138) );
  OAI221XL U193 ( .A0(n5203), .A1(n4783), .B0(n5202), .B1(n5007), .C0(n1142), 
        .Y(n1137) );
  OAI221XL U194 ( .A0(n5219), .A1(n4784), .B0(n5218), .B1(n5008), .C0(n1140), 
        .Y(n1139) );
  OR4X2 U195 ( .A(n1128), .B(n1129), .C(n1130), .D(n1131), .Y(\rd2<26> ) );
  OAI221XL U196 ( .A0(n5211), .A1(n4785), .B0(n5210), .B1(n5009), .C0(n1133), 
        .Y(n1130) );
  OAI221XL U197 ( .A0(n5203), .A1(n4786), .B0(n5202), .B1(n5010), .C0(n1134), 
        .Y(n1129) );
  OAI221XL U198 ( .A0(n5219), .A1(n4787), .B0(n5218), .B1(n5011), .C0(n1132), 
        .Y(n1131) );
  BUFX3 U199 ( .A(\wd3<18> ), .Y(n5128) );
  BUFX3 U200 ( .A(\wd3<19> ), .Y(n5129) );
  BUFX3 U201 ( .A(\wd3<20> ), .Y(n5130) );
  BUFX3 U202 ( .A(\wd3<21> ), .Y(n5131) );
  BUFX3 U203 ( .A(\wd3<22> ), .Y(n5132) );
  OR4X2 U204 ( .A(n1208), .B(n1209), .C(n1210), .D(n1211), .Y(\rd2<17> ) );
  OAI221XL U205 ( .A0(n5212), .A1(n4788), .B0(n5209), .B1(n5012), .C0(n1213), 
        .Y(n1210) );
  OAI221XL U206 ( .A0(n5204), .A1(n4789), .B0(n5201), .B1(n5013), .C0(n1214), 
        .Y(n1209) );
  OAI221XL U207 ( .A0(n5220), .A1(n4790), .B0(n5217), .B1(n5014), .C0(n1212), 
        .Y(n1211) );
  OR4X2 U208 ( .A(n1200), .B(n1201), .C(n1202), .D(n1203), .Y(\rd2<18> ) );
  OAI221XL U209 ( .A0(n5212), .A1(n4791), .B0(n5209), .B1(n5015), .C0(n1205), 
        .Y(n1202) );
  OAI221XL U210 ( .A0(n5204), .A1(n4792), .B0(n5201), .B1(n5016), .C0(n1206), 
        .Y(n1201) );
  OAI221XL U211 ( .A0(n5220), .A1(n4793), .B0(n5217), .B1(n5017), .C0(n1204), 
        .Y(n1203) );
  OR4X2 U212 ( .A(n1192), .B(n1193), .C(n1194), .D(n1195), .Y(\rd2<19> ) );
  OAI221XL U213 ( .A0(n5212), .A1(n4794), .B0(n5209), .B1(n5018), .C0(n1197), 
        .Y(n1194) );
  OAI221XL U214 ( .A0(n5204), .A1(n4795), .B0(n5201), .B1(n5019), .C0(n1198), 
        .Y(n1193) );
  OAI221XL U215 ( .A0(n5220), .A1(n4796), .B0(n5217), .B1(n5020), .C0(n1196), 
        .Y(n1195) );
  OR4X2 U216 ( .A(n1176), .B(n1177), .C(n1178), .D(n1179), .Y(\rd2<20> ) );
  OAI221XL U217 ( .A0(n5211), .A1(n4797), .B0(n5210), .B1(n5021), .C0(n1181), 
        .Y(n1178) );
  OAI221XL U218 ( .A0(n5203), .A1(n4798), .B0(n5202), .B1(n5022), .C0(n1182), 
        .Y(n1177) );
  OAI221XL U219 ( .A0(n5219), .A1(n4799), .B0(n5218), .B1(n5023), .C0(n1180), 
        .Y(n1179) );
  OR4X2 U220 ( .A(n1168), .B(n1169), .C(n1170), .D(n1171), .Y(\rd2<21> ) );
  OAI221XL U221 ( .A0(n5211), .A1(n4800), .B0(n5210), .B1(n5024), .C0(n1173), 
        .Y(n1170) );
  OAI221XL U222 ( .A0(n5203), .A1(n4801), .B0(n5202), .B1(n5025), .C0(n1174), 
        .Y(n1169) );
  OAI221XL U223 ( .A0(n5219), .A1(n4802), .B0(n5218), .B1(n5026), .C0(n1172), 
        .Y(n1171) );
  BUFX3 U224 ( .A(\wd3<13> ), .Y(n5123) );
  BUFX3 U225 ( .A(\wd3<14> ), .Y(n5124) );
  BUFX3 U226 ( .A(\wd3<15> ), .Y(n5125) );
  BUFX3 U227 ( .A(\wd3<16> ), .Y(n5126) );
  BUFX3 U228 ( .A(\wd3<17> ), .Y(n5127) );
  OR4X2 U229 ( .A(n1248), .B(n1249), .C(n1250), .D(n1251), .Y(\rd2<12> ) );
  OAI221XL U230 ( .A0(n5212), .A1(n4803), .B0(n5209), .B1(n5027), .C0(n1253), 
        .Y(n1250) );
  OAI221XL U231 ( .A0(n5204), .A1(n4804), .B0(n5201), .B1(n5028), .C0(n1254), 
        .Y(n1249) );
  OAI221XL U232 ( .A0(n5220), .A1(n4805), .B0(n5217), .B1(n5029), .C0(n1252), 
        .Y(n1251) );
  OR4X2 U233 ( .A(n1240), .B(n1241), .C(n1242), .D(n1243), .Y(\rd2<13> ) );
  OAI221XL U234 ( .A0(n5211), .A1(n4806), .B0(n5209), .B1(n5030), .C0(n1245), 
        .Y(n1242) );
  OAI221XL U235 ( .A0(n5203), .A1(n4807), .B0(n5201), .B1(n5031), .C0(n1246), 
        .Y(n1241) );
  OAI221XL U236 ( .A0(n5219), .A1(n4808), .B0(n5217), .B1(n5032), .C0(n1244), 
        .Y(n1243) );
  OR4X2 U237 ( .A(n1232), .B(n1233), .C(n1234), .D(n1235), .Y(\rd2<14> ) );
  OAI221XL U238 ( .A0(n5212), .A1(n4809), .B0(n5209), .B1(n5033), .C0(n1237), 
        .Y(n1234) );
  OAI221XL U239 ( .A0(n5204), .A1(n4810), .B0(n5201), .B1(n5034), .C0(n1238), 
        .Y(n1233) );
  OAI221XL U240 ( .A0(n5220), .A1(n4811), .B0(n5217), .B1(n5035), .C0(n1236), 
        .Y(n1235) );
  OR4X2 U241 ( .A(n1224), .B(n1225), .C(n1226), .D(n1227), .Y(\rd2<15> ) );
  OAI221XL U242 ( .A0(n5211), .A1(n4812), .B0(n5209), .B1(n5036), .C0(n1229), 
        .Y(n1226) );
  OAI221XL U243 ( .A0(n5203), .A1(n4813), .B0(n5201), .B1(n5037), .C0(n1230), 
        .Y(n1225) );
  OAI221XL U244 ( .A0(n5219), .A1(n4814), .B0(n5217), .B1(n5038), .C0(n1228), 
        .Y(n1227) );
  OR4X2 U245 ( .A(n1216), .B(n1217), .C(n1218), .D(n1219), .Y(\rd2<16> ) );
  OAI221XL U246 ( .A0(n5212), .A1(n4815), .B0(n5209), .B1(n5039), .C0(n1221), 
        .Y(n1218) );
  OAI221XL U247 ( .A0(n5204), .A1(n4816), .B0(n5201), .B1(n5040), .C0(n1222), 
        .Y(n1217) );
  OAI221XL U248 ( .A0(n5220), .A1(n4817), .B0(n5217), .B1(n5041), .C0(n1220), 
        .Y(n1219) );
  BUFX3 U249 ( .A(\wd3<7> ), .Y(n5117) );
  BUFX3 U250 ( .A(\wd3<8> ), .Y(n5118) );
  BUFX3 U251 ( .A(\wd3<9> ), .Y(n5119) );
  BUFX3 U252 ( .A(\wd3<10> ), .Y(n5120) );
  BUFX3 U253 ( .A(\wd3<11> ), .Y(n5121) );
  BUFX3 U254 ( .A(\wd3<12> ), .Y(n5122) );
  OR4X2 U255 ( .A(n1048), .B(n1049), .C(n1050), .D(n1051), .Y(\rd2<6> ) );
  OAI221XL U256 ( .A0(n5212), .A1(n4818), .B0(n5209), .B1(n5042), .C0(n1053), 
        .Y(n1050) );
  OAI221XL U257 ( .A0(n5204), .A1(n4819), .B0(n5201), .B1(n5043), .C0(n1054), 
        .Y(n1049) );
  OAI221XL U258 ( .A0(n5220), .A1(n4820), .B0(n5217), .B1(n5044), .C0(n1052), 
        .Y(n1051) );
  OR4X2 U259 ( .A(n1040), .B(n1041), .C(n1042), .D(n1043), .Y(\rd2<7> ) );
  OAI221XL U260 ( .A0(n5212), .A1(n4821), .B0(n5210), .B1(n5045), .C0(n1045), 
        .Y(n1042) );
  OAI221XL U261 ( .A0(n5204), .A1(n4822), .B0(n5202), .B1(n5046), .C0(n1046), 
        .Y(n1041) );
  OAI221XL U262 ( .A0(n5220), .A1(n4823), .B0(n5218), .B1(n5047), .C0(n1044), 
        .Y(n1043) );
  OR4X2 U263 ( .A(n1032), .B(n1033), .C(n1034), .D(n1035), .Y(\rd2<8> ) );
  OAI221XL U264 ( .A0(n5212), .A1(n4824), .B0(n5209), .B1(n5048), .C0(n1037), 
        .Y(n1034) );
  OAI221XL U265 ( .A0(n5204), .A1(n4825), .B0(n5201), .B1(n5049), .C0(n1038), 
        .Y(n1033) );
  OAI221XL U266 ( .A0(n5220), .A1(n4826), .B0(n5217), .B1(n5050), .C0(n1036), 
        .Y(n1035) );
  OR4X2 U267 ( .A(n1008), .B(n1009), .C(n1010), .D(n1011), .Y(\rd2<9> ) );
  OAI221XL U268 ( .A0(n5212), .A1(n4827), .B0(n5210), .B1(n5051), .C0(n1019), 
        .Y(n1010) );
  OAI221XL U269 ( .A0(n5204), .A1(n4828), .B0(n5202), .B1(n5052), .C0(n1024), 
        .Y(n1009) );
  OAI221XL U270 ( .A0(n5220), .A1(n4829), .B0(n5218), .B1(n5053), .C0(n1014), 
        .Y(n1011) );
  OR4X2 U271 ( .A(n1264), .B(n1265), .C(n1266), .D(n1267), .Y(\rd2<10> ) );
  OAI221XL U272 ( .A0(n5211), .A1(n4830), .B0(n5209), .B1(n5054), .C0(n1269), 
        .Y(n1266) );
  OAI221XL U273 ( .A0(n5203), .A1(n4831), .B0(n5201), .B1(n5055), .C0(n1270), 
        .Y(n1265) );
  OAI221XL U274 ( .A0(n5219), .A1(n4832), .B0(n5217), .B1(n5056), .C0(n1268), 
        .Y(n1267) );
  OR4X2 U275 ( .A(n1256), .B(n1257), .C(n1258), .D(n1259), .Y(\rd2<11> ) );
  OAI221XL U276 ( .A0(n5212), .A1(n4833), .B0(n5209), .B1(n5057), .C0(n1261), 
        .Y(n1258) );
  OAI221XL U277 ( .A0(n5204), .A1(n4834), .B0(n5201), .B1(n5058), .C0(n1262), 
        .Y(n1257) );
  OAI221XL U278 ( .A0(n5220), .A1(n4835), .B0(n5217), .B1(n5059), .C0(n1260), 
        .Y(n1259) );
  BUFX3 U279 ( .A(\wd3<2> ), .Y(n5112) );
  BUFX3 U280 ( .A(\wd3<3> ), .Y(n5113) );
  BUFX3 U281 ( .A(\wd3<4> ), .Y(n5114) );
  BUFX3 U282 ( .A(\wd3<5> ), .Y(n5115) );
  BUFX3 U283 ( .A(\wd3<6> ), .Y(n5116) );
  OR4X2 U284 ( .A(n1184), .B(n1185), .C(n1186), .D(n1187), .Y(\rd2<1> ) );
  OAI221XL U285 ( .A0(n5211), .A1(n4836), .B0(n5209), .B1(n5060), .C0(n1189), 
        .Y(n1186) );
  OAI221XL U286 ( .A0(n5203), .A1(n4837), .B0(n5201), .B1(n5061), .C0(n1190), 
        .Y(n1185) );
  OAI221XL U287 ( .A0(n5219), .A1(n4838), .B0(n5217), .B1(n5062), .C0(n1188), 
        .Y(n1187) );
  OR4X2 U288 ( .A(n1096), .B(n1097), .C(n1098), .D(n1099), .Y(\rd2<2> ) );
  OAI221XL U289 ( .A0(n5211), .A1(n4839), .B0(n5210), .B1(n5063), .C0(n1101), 
        .Y(n1098) );
  OAI221XL U290 ( .A0(n5203), .A1(n4840), .B0(n5202), .B1(n5064), .C0(n1102), 
        .Y(n1097) );
  OAI221XL U291 ( .A0(n5219), .A1(n4841), .B0(n5218), .B1(n5065), .C0(n1100), 
        .Y(n1099) );
  OR4X2 U292 ( .A(n1072), .B(n1073), .C(n1074), .D(n1075), .Y(\rd2<3> ) );
  OAI221XL U293 ( .A0(n5212), .A1(n4842), .B0(n5209), .B1(n5066), .C0(n1077), 
        .Y(n1074) );
  OAI221XL U294 ( .A0(n5204), .A1(n4843), .B0(n5201), .B1(n5067), .C0(n1078), 
        .Y(n1073) );
  OAI221XL U295 ( .A0(n5220), .A1(n4844), .B0(n5217), .B1(n5068), .C0(n1076), 
        .Y(n1075) );
  OR4X2 U296 ( .A(n1064), .B(n1065), .C(n1066), .D(n1067), .Y(\rd2<4> ) );
  OAI221XL U297 ( .A0(n5212), .A1(n4845), .B0(n5210), .B1(n5069), .C0(n1069), 
        .Y(n1066) );
  OAI221XL U298 ( .A0(n5204), .A1(n4846), .B0(n5202), .B1(n5070), .C0(n1070), 
        .Y(n1065) );
  OAI221XL U299 ( .A0(n5220), .A1(n4847), .B0(n5218), .B1(n5071), .C0(n1068), 
        .Y(n1067) );
  OR4X2 U300 ( .A(n1056), .B(n1057), .C(n1058), .D(n1059), .Y(\rd2<5> ) );
  OAI221XL U301 ( .A0(n5212), .A1(n4848), .B0(n5209), .B1(n5072), .C0(n1061), 
        .Y(n1058) );
  OAI221XL U302 ( .A0(n5204), .A1(n4849), .B0(n5201), .B1(n5073), .C0(n1062), 
        .Y(n1057) );
  OAI221XL U303 ( .A0(n5220), .A1(n4850), .B0(n5217), .B1(n5074), .C0(n1060), 
        .Y(n1059) );
  BUFX3 U304 ( .A(\wd3<0> ), .Y(n5110) );
  BUFX3 U305 ( .A(\wd3<1> ), .Y(n5111) );
  OR4X2 U306 ( .A(n1272), .B(n1273), .C(n1274), .D(n1275), .Y(\rd2<0> ) );
  OAI221XL U307 ( .A0(n5212), .A1(n4851), .B0(n5209), .B1(n5075), .C0(n1280), 
        .Y(n1274) );
  OAI221XL U308 ( .A0(n5204), .A1(n4852), .B0(n5201), .B1(n5076), .C0(n1282), 
        .Y(n1273) );
  OAI221XL U309 ( .A0(n5220), .A1(n4853), .B0(n5217), .B1(n5077), .C0(n1276), 
        .Y(n1275) );
  NOR2X1 U310 ( .A(N12), .B(N13), .Y(n1557) );
  NOR2X1 U311 ( .A(n5282), .B(N13), .Y(n1558) );
  NOR2X1 U312 ( .A(n5290), .B(N18), .Y(n1279) );
  NAND3X1 U313 ( .A(n5287), .B(n5285), .C(we3), .Y(n1564) );
  NOR2X1 U314 ( .A(n5280), .B(N14), .Y(n1562) );
  NOR2X1 U315 ( .A(n5281), .B(N15), .Y(n1560) );
  NOR2X1 U316 ( .A(N14), .B(N15), .Y(n1555) );
  NOR2X1 U317 ( .A(n5284), .B(N19), .Y(n1281) );
  NOR3X1 U318 ( .A(n5284), .B(N17), .C(n5286), .Y(n1277) );
  CLKINVX3 U319 ( .A(n5142), .Y(n5288) );
  CLKINVX3 U320 ( .A(N17), .Y(n5290) );
  AND2X2 U321 ( .A(N13), .B(N12), .Y(n1556) );
  AND2X2 U322 ( .A(N13), .B(n5282), .Y(n1554) );
  NOR2X1 U323 ( .A(n1568), .B(n1571), .Y(n1580) );
  NOR2X1 U324 ( .A(n1565), .B(n1568), .Y(n15) );
  NOR2X1 U325 ( .A(n1566), .B(n1568), .Y(n1575) );
  NOR2X1 U326 ( .A(n1567), .B(n1568), .Y(n1579) );
  NOR2X1 U327 ( .A(n1565), .B(n1569), .Y(n16) );
  NOR2X1 U328 ( .A(n1564), .B(n1567), .Y(n1574) );
  NOR2X1 U329 ( .A(n1564), .B(n1565), .Y(n1572) );
  NOR2X1 U330 ( .A(n1564), .B(n1571), .Y(n13) );
  INVX1 U331 ( .A(N19), .Y(n5286) );
  NAND3X1 U332 ( .A(n1279), .B(n5288), .C(N19), .Y(n1028) );
  INVX1 U333 ( .A(N15), .Y(n5280) );
  INVX1 U334 ( .A(N14), .Y(n5281) );
  INVX1 U335 ( .A(N12), .Y(n5282) );
  NAND2X1 U336 ( .A(n5289), .B(n5283), .Y(n1566) );
  OAI221XL U337 ( .A0(n4099), .A1(n5163), .B0(n3939), .B1(n5159), .C0(n1363), 
        .Y(n1356) );
  AOI22X1 U338 ( .A0(n5157), .A1(\r15<31> ), .B0(n1307), .B1(\rf<10><31> ), 
        .Y(n1363) );
  OAI221XL U339 ( .A0(n5196), .A1(n5248), .B0(n5193), .B1(n5078), .C0(n1087), 
        .Y(n1080) );
  AOI22X1 U340 ( .A0(n5191), .A1(n4630), .B0(n5189), .B1(n4854), .Y(n1087) );
  INVX1 U341 ( .A(\r15<31> ), .Y(n5248) );
  OR4X2 U342 ( .A(n1356), .B(n1357), .C(n1358), .D(n1359), .Y(\rd1<31> ) );
  OAI221XL U343 ( .A0(n4100), .A1(n5171), .B0(n3940), .B1(n5169), .C0(n1362), 
        .Y(n1357) );
  OAI221XL U344 ( .A0(n4101), .A1(n5179), .B0(n3941), .B1(n5177), .C0(n1361), 
        .Y(n1358) );
  OAI221XL U345 ( .A0(n4354), .A1(n5187), .B0(n4322), .B1(n5185), .C0(n1360), 
        .Y(n1359) );
  OAI221XL U346 ( .A0(n4107), .A1(n5163), .B0(n3947), .B1(n5159), .C0(n1403), 
        .Y(n1396) );
  AOI22X1 U347 ( .A0(n5157), .A1(\r15<27> ), .B0(n5155), .B1(\rf<10><27> ), 
        .Y(n1403) );
  OAI221XL U348 ( .A0(n4108), .A1(n5163), .B0(n3948), .B1(n5159), .C0(n1395), 
        .Y(n1388) );
  AOI22X1 U349 ( .A0(n5157), .A1(\r15<28> ), .B0(n5155), .B1(\rf<10><28> ), 
        .Y(n1395) );
  OAI221XL U350 ( .A0(n4109), .A1(n5163), .B0(n3949), .B1(n5159), .C0(n1387), 
        .Y(n1380) );
  AOI22X1 U351 ( .A0(n5157), .A1(\r15<29> ), .B0(n5155), .B1(\rf<10><29> ), 
        .Y(n1387) );
  OAI221XL U352 ( .A0(n4102), .A1(n5163), .B0(n3942), .B1(n5159), .C0(n1371), 
        .Y(n1364) );
  AOI22X1 U353 ( .A0(n5157), .A1(\r15<30> ), .B0(n5155), .B1(\rf<10><30> ), 
        .Y(n1371) );
  OAI221XL U354 ( .A0(n5196), .A1(n5252), .B0(n5193), .B1(n5079), .C0(n1127), 
        .Y(n1120) );
  AOI22X1 U355 ( .A0(n5190), .A1(n4631), .B0(n5189), .B1(n4855), .Y(n1127) );
  INVX1 U356 ( .A(\r15<27> ), .Y(n5252) );
  OAI221XL U357 ( .A0(n5196), .A1(n5251), .B0(n5193), .B1(n5080), .C0(n1119), 
        .Y(n1112) );
  AOI22X1 U358 ( .A0(n5190), .A1(n4632), .B0(n5189), .B1(n4856), .Y(n1119) );
  INVX1 U359 ( .A(\r15<28> ), .Y(n5251) );
  OAI221XL U360 ( .A0(n5196), .A1(n5250), .B0(n5193), .B1(n5081), .C0(n1111), 
        .Y(n1104) );
  AOI22X1 U361 ( .A0(n5190), .A1(n4633), .B0(n5189), .B1(n4857), .Y(n1111) );
  INVX1 U362 ( .A(\r15<29> ), .Y(n5250) );
  OAI221XL U363 ( .A0(n5196), .A1(n5249), .B0(n5193), .B1(n5082), .C0(n1095), 
        .Y(n1088) );
  AOI22X1 U364 ( .A0(n5190), .A1(n4634), .B0(n5189), .B1(n4858), .Y(n1095) );
  INVX1 U365 ( .A(\r15<30> ), .Y(n5249) );
  OR4X2 U366 ( .A(n1396), .B(n1397), .C(n1398), .D(n1399), .Y(\rd1<27> ) );
  OAI221XL U367 ( .A0(n4114), .A1(n5171), .B0(n3954), .B1(n5169), .C0(n1402), 
        .Y(n1397) );
  OAI221XL U368 ( .A0(n4115), .A1(n5179), .B0(n3955), .B1(n5177), .C0(n1401), 
        .Y(n1398) );
  OAI221XL U369 ( .A0(n4350), .A1(n5187), .B0(n4318), .B1(n5185), .C0(n1400), 
        .Y(n1399) );
  OR4X2 U370 ( .A(n1388), .B(n1389), .C(n1390), .D(n1391), .Y(\rd1<28> ) );
  OAI221XL U371 ( .A0(n4116), .A1(n5171), .B0(n3956), .B1(n5169), .C0(n1394), 
        .Y(n1389) );
  OAI221XL U372 ( .A0(n4117), .A1(n5179), .B0(n3957), .B1(n5177), .C0(n1393), 
        .Y(n1390) );
  OAI221XL U373 ( .A0(n4351), .A1(n5187), .B0(n4319), .B1(n5185), .C0(n1392), 
        .Y(n1391) );
  OR4X2 U374 ( .A(n1380), .B(n1381), .C(n1382), .D(n1383), .Y(\rd1<29> ) );
  OAI221XL U375 ( .A0(n4118), .A1(n5171), .B0(n3958), .B1(n5169), .C0(n1386), 
        .Y(n1381) );
  OAI221XL U376 ( .A0(n4119), .A1(n5179), .B0(n3959), .B1(n5177), .C0(n1385), 
        .Y(n1382) );
  OAI221XL U377 ( .A0(n4352), .A1(n5187), .B0(n4320), .B1(n5185), .C0(n1384), 
        .Y(n1383) );
  OR4X2 U378 ( .A(n1364), .B(n1365), .C(n1366), .D(n1367), .Y(\rd1<30> ) );
  OAI221XL U379 ( .A0(n4103), .A1(n5171), .B0(n3943), .B1(n5169), .C0(n1370), 
        .Y(n1365) );
  OAI221XL U380 ( .A0(n4104), .A1(n5179), .B0(n3944), .B1(n5177), .C0(n1369), 
        .Y(n1366) );
  OAI221XL U381 ( .A0(n4353), .A1(n5187), .B0(n4321), .B1(n5185), .C0(n1368), 
        .Y(n1367) );
  OAI221XL U382 ( .A0(n4122), .A1(n5163), .B0(n3962), .B1(n5159), .C0(n1443), 
        .Y(n1436) );
  AOI22X1 U383 ( .A0(n5157), .A1(\r15<22> ), .B0(n5155), .B1(\rf<10><22> ), 
        .Y(n1443) );
  OAI221XL U384 ( .A0(n4123), .A1(n5163), .B0(n3963), .B1(n5159), .C0(n1435), 
        .Y(n1428) );
  AOI22X1 U385 ( .A0(n5157), .A1(\r15<23> ), .B0(n5155), .B1(\rf<10><23> ), 
        .Y(n1435) );
  OAI221XL U386 ( .A0(n4124), .A1(n5163), .B0(n3964), .B1(n5159), .C0(n1427), 
        .Y(n1420) );
  AOI22X1 U387 ( .A0(n5157), .A1(\r15<24> ), .B0(n5155), .B1(\rf<10><24> ), 
        .Y(n1427) );
  OAI221XL U388 ( .A0(n4105), .A1(n5163), .B0(n3945), .B1(n5159), .C0(n1419), 
        .Y(n1412) );
  AOI22X1 U389 ( .A0(n5157), .A1(\r15<25> ), .B0(n5155), .B1(\rf<10><25> ), 
        .Y(n1419) );
  OAI221XL U390 ( .A0(n4106), .A1(n5163), .B0(n3946), .B1(n5159), .C0(n1411), 
        .Y(n1404) );
  AOI22X1 U391 ( .A0(n5157), .A1(\r15<26> ), .B0(n5155), .B1(\rf<10><26> ), 
        .Y(n1411) );
  OAI221XL U392 ( .A0(n5196), .A1(n5257), .B0(n5193), .B1(n5083), .C0(n1167), 
        .Y(n1160) );
  AOI22X1 U393 ( .A0(n5190), .A1(n4635), .B0(n5189), .B1(n4859), .Y(n1167) );
  INVX1 U394 ( .A(\r15<22> ), .Y(n5257) );
  OAI221XL U395 ( .A0(n5196), .A1(n5256), .B0(n5193), .B1(n5084), .C0(n1159), 
        .Y(n1152) );
  AOI22X1 U396 ( .A0(n5190), .A1(n4636), .B0(n5189), .B1(n4860), .Y(n1159) );
  INVX1 U397 ( .A(\r15<23> ), .Y(n5256) );
  OAI221XL U398 ( .A0(n5196), .A1(n5255), .B0(n5193), .B1(n5085), .C0(n1151), 
        .Y(n1144) );
  AOI22X1 U399 ( .A0(n5190), .A1(n4637), .B0(n5189), .B1(n4861), .Y(n1151) );
  INVX1 U400 ( .A(\r15<24> ), .Y(n5255) );
  OAI221XL U401 ( .A0(n5196), .A1(n5254), .B0(n5193), .B1(n5086), .C0(n1143), 
        .Y(n1136) );
  AOI22X1 U402 ( .A0(n5190), .A1(n4638), .B0(n5189), .B1(n4862), .Y(n1143) );
  INVX1 U403 ( .A(\r15<25> ), .Y(n5254) );
  OAI221XL U404 ( .A0(n5196), .A1(n5253), .B0(n5193), .B1(n5087), .C0(n1135), 
        .Y(n1128) );
  AOI22X1 U405 ( .A0(n5190), .A1(n4639), .B0(n5189), .B1(n4863), .Y(n1135) );
  INVX1 U406 ( .A(\r15<26> ), .Y(n5253) );
  OR4X2 U407 ( .A(n1436), .B(n1437), .C(n1438), .D(n1439), .Y(\rd1<22> ) );
  OAI221XL U408 ( .A0(n4129), .A1(n5171), .B0(n3969), .B1(n5169), .C0(n1442), 
        .Y(n1437) );
  OAI221XL U409 ( .A0(n4130), .A1(n5179), .B0(n3970), .B1(n5177), .C0(n1441), 
        .Y(n1438) );
  OAI221XL U410 ( .A0(n4345), .A1(n5187), .B0(n4313), .B1(n5185), .C0(n1440), 
        .Y(n1439) );
  OR4X2 U411 ( .A(n1428), .B(n1429), .C(n1430), .D(n1431), .Y(\rd1<23> ) );
  OAI221XL U412 ( .A0(n4131), .A1(n5171), .B0(n3971), .B1(n5169), .C0(n1434), 
        .Y(n1429) );
  OAI221XL U413 ( .A0(n4132), .A1(n5179), .B0(n3972), .B1(n5177), .C0(n1433), 
        .Y(n1430) );
  OAI221XL U414 ( .A0(n4346), .A1(n5187), .B0(n4314), .B1(n5185), .C0(n1432), 
        .Y(n1431) );
  OR4X2 U415 ( .A(n1420), .B(n1421), .C(n1422), .D(n1423), .Y(\rd1<24> ) );
  OAI221XL U416 ( .A0(n4133), .A1(n5171), .B0(n3973), .B1(n5169), .C0(n1426), 
        .Y(n1421) );
  OAI221XL U417 ( .A0(n4134), .A1(n5179), .B0(n3974), .B1(n5177), .C0(n1425), 
        .Y(n1422) );
  OAI221XL U418 ( .A0(n4347), .A1(n5187), .B0(n4315), .B1(n5185), .C0(n1424), 
        .Y(n1423) );
  OR4X2 U419 ( .A(n1412), .B(n1413), .C(n1414), .D(n1415), .Y(\rd1<25> ) );
  OAI221XL U420 ( .A0(n4110), .A1(n5171), .B0(n3950), .B1(n5169), .C0(n1418), 
        .Y(n1413) );
  OAI221XL U421 ( .A0(n4111), .A1(n5179), .B0(n3951), .B1(n5177), .C0(n1417), 
        .Y(n1414) );
  OAI221XL U422 ( .A0(n4348), .A1(n5187), .B0(n4316), .B1(n5185), .C0(n1416), 
        .Y(n1415) );
  OR4X2 U423 ( .A(n1404), .B(n1405), .C(n1406), .D(n1407), .Y(\rd1<26> ) );
  OAI221XL U424 ( .A0(n4112), .A1(n5171), .B0(n3952), .B1(n5169), .C0(n1410), 
        .Y(n1405) );
  OAI221XL U425 ( .A0(n4113), .A1(n5179), .B0(n3953), .B1(n5177), .C0(n1409), 
        .Y(n1406) );
  OAI221XL U426 ( .A0(n4349), .A1(n5187), .B0(n4317), .B1(n5185), .C0(n1408), 
        .Y(n1407) );
  OAI221XL U427 ( .A0(n4136), .A1(n5162), .B0(n3976), .B1(n5160), .C0(n1499), 
        .Y(n1492) );
  AOI22X1 U428 ( .A0(n5157), .A1(\r15<16> ), .B0(n1307), .B1(\rf<10><16> ), 
        .Y(n1499) );
  OAI221XL U429 ( .A0(n4137), .A1(n5162), .B0(n3977), .B1(n5159), .C0(n1491), 
        .Y(n1484) );
  AOI22X1 U430 ( .A0(n5157), .A1(\r15<17> ), .B0(n1307), .B1(\rf<10><17> ), 
        .Y(n1491) );
  OAI221XL U431 ( .A0(n4138), .A1(n5162), .B0(n3978), .B1(n5159), .C0(n1483), 
        .Y(n1476) );
  AOI22X1 U432 ( .A0(n5157), .A1(\r15<18> ), .B0(n1307), .B1(\rf<10><18> ), 
        .Y(n1483) );
  OAI221XL U433 ( .A0(n4139), .A1(n5162), .B0(n3979), .B1(n5159), .C0(n1475), 
        .Y(n1468) );
  AOI22X1 U434 ( .A0(n5157), .A1(\r15<19> ), .B0(n1307), .B1(\rf<10><19> ), 
        .Y(n1475) );
  OAI221XL U435 ( .A0(n4120), .A1(n5162), .B0(n3960), .B1(n1304), .C0(n1459), 
        .Y(n1452) );
  AOI22X1 U436 ( .A0(n5157), .A1(\r15<20> ), .B0(n5155), .B1(\rf<10><20> ), 
        .Y(n1459) );
  OAI221XL U437 ( .A0(n4121), .A1(n5163), .B0(n3961), .B1(n5159), .C0(n1451), 
        .Y(n1444) );
  AOI22X1 U438 ( .A0(n5157), .A1(\r15<21> ), .B0(n5155), .B1(\rf<10><21> ), 
        .Y(n1451) );
  OAI221XL U439 ( .A0(n5195), .A1(n5262), .B0(n5192), .B1(n5088), .C0(n1215), 
        .Y(n1208) );
  AOI22X1 U440 ( .A0(n5191), .A1(n4640), .B0(n5188), .B1(n4864), .Y(n1215) );
  INVX1 U441 ( .A(\r15<17> ), .Y(n5262) );
  OAI221XL U442 ( .A0(n5195), .A1(n5261), .B0(n5192), .B1(n5089), .C0(n1207), 
        .Y(n1200) );
  AOI22X1 U443 ( .A0(n5191), .A1(n4641), .B0(n5188), .B1(n4865), .Y(n1207) );
  INVX1 U444 ( .A(\r15<18> ), .Y(n5261) );
  OAI221XL U445 ( .A0(n5195), .A1(n5260), .B0(n5192), .B1(n5090), .C0(n1199), 
        .Y(n1192) );
  AOI22X1 U446 ( .A0(n5191), .A1(n4642), .B0(n5188), .B1(n4866), .Y(n1199) );
  INVX1 U447 ( .A(\r15<19> ), .Y(n5260) );
  OAI221XL U448 ( .A0(n5196), .A1(n5259), .B0(n5193), .B1(n5091), .C0(n1183), 
        .Y(n1176) );
  AOI22X1 U449 ( .A0(n5190), .A1(n4643), .B0(n5189), .B1(n4867), .Y(n1183) );
  INVX1 U450 ( .A(\r15<20> ), .Y(n5259) );
  OAI221XL U451 ( .A0(n5196), .A1(n5258), .B0(n5193), .B1(n5092), .C0(n1175), 
        .Y(n1168) );
  AOI22X1 U452 ( .A0(n5190), .A1(n4644), .B0(n5189), .B1(n4868), .Y(n1175) );
  INVX1 U453 ( .A(\r15<21> ), .Y(n5258) );
  OR4X2 U454 ( .A(n1492), .B(n1493), .C(n1494), .D(n1495), .Y(\rd1<16> ) );
  OAI221XL U455 ( .A0(n4142), .A1(n5170), .B0(n3982), .B1(n5168), .C0(n1498), 
        .Y(n1493) );
  OAI221XL U456 ( .A0(n4143), .A1(n5178), .B0(n3983), .B1(n5176), .C0(n1497), 
        .Y(n1494) );
  OAI221XL U457 ( .A0(n4339), .A1(n5186), .B0(n4307), .B1(n5184), .C0(n1496), 
        .Y(n1495) );
  OR4X2 U458 ( .A(n1484), .B(n1485), .C(n1486), .D(n1487), .Y(\rd1<17> ) );
  OAI221XL U459 ( .A0(n4144), .A1(n5170), .B0(n3984), .B1(n5168), .C0(n1490), 
        .Y(n1485) );
  OAI221XL U460 ( .A0(n4145), .A1(n5178), .B0(n3985), .B1(n5176), .C0(n1489), 
        .Y(n1486) );
  OAI221XL U461 ( .A0(n4340), .A1(n5186), .B0(n4308), .B1(n5184), .C0(n1488), 
        .Y(n1487) );
  OR4X2 U462 ( .A(n1476), .B(n1477), .C(n1478), .D(n1479), .Y(\rd1<18> ) );
  OAI221XL U463 ( .A0(n4146), .A1(n5170), .B0(n3986), .B1(n5168), .C0(n1482), 
        .Y(n1477) );
  OAI221XL U464 ( .A0(n4147), .A1(n5178), .B0(n3987), .B1(n5176), .C0(n1481), 
        .Y(n1478) );
  OAI221XL U465 ( .A0(n4341), .A1(n5186), .B0(n4309), .B1(n5184), .C0(n1480), 
        .Y(n1479) );
  OR4X2 U466 ( .A(n1468), .B(n1469), .C(n1470), .D(n1471), .Y(\rd1<19> ) );
  OAI221XL U467 ( .A0(n4148), .A1(n5170), .B0(n3988), .B1(n5168), .C0(n1474), 
        .Y(n1469) );
  OAI221XL U468 ( .A0(n4149), .A1(n5178), .B0(n3989), .B1(n5176), .C0(n1473), 
        .Y(n1470) );
  OAI221XL U469 ( .A0(n4342), .A1(n5186), .B0(n4310), .B1(n5184), .C0(n1472), 
        .Y(n1471) );
  OR4X2 U470 ( .A(n1452), .B(n1453), .C(n1454), .D(n1455), .Y(\rd1<20> ) );
  OAI221XL U471 ( .A0(n4125), .A1(n5170), .B0(n3965), .B1(n5168), .C0(n1458), 
        .Y(n1453) );
  OAI221XL U472 ( .A0(n4126), .A1(n5178), .B0(n3966), .B1(n5176), .C0(n1457), 
        .Y(n1454) );
  OAI221XL U473 ( .A0(n4343), .A1(n5186), .B0(n4311), .B1(n5184), .C0(n1456), 
        .Y(n1455) );
  OR4X2 U474 ( .A(n1444), .B(n1445), .C(n1446), .D(n1447), .Y(\rd1<21> ) );
  OAI221XL U475 ( .A0(n4127), .A1(n5171), .B0(n3967), .B1(n5169), .C0(n1450), 
        .Y(n1445) );
  OAI221XL U476 ( .A0(n4128), .A1(n5179), .B0(n3968), .B1(n5177), .C0(n1449), 
        .Y(n1446) );
  OAI221XL U477 ( .A0(n4344), .A1(n5187), .B0(n4312), .B1(n5185), .C0(n1448), 
        .Y(n1447) );
  OAI221XL U478 ( .A0(n4151), .A1(n5162), .B0(n3991), .B1(n1304), .C0(n1539), 
        .Y(n1532) );
  AOI22X1 U479 ( .A0(n1306), .A1(\r15<11> ), .B0(n5155), .B1(\rf<10><11> ), 
        .Y(n1539) );
  OAI221XL U480 ( .A0(n4152), .A1(n5162), .B0(n3992), .B1(n1304), .C0(n1531), 
        .Y(n1524) );
  AOI22X1 U481 ( .A0(n1306), .A1(\r15<12> ), .B0(n5155), .B1(\rf<10><12> ), 
        .Y(n1531) );
  OAI221XL U482 ( .A0(n4153), .A1(n5162), .B0(n3993), .B1(n1304), .C0(n1523), 
        .Y(n1516) );
  AOI22X1 U483 ( .A0(n1306), .A1(\r15<13> ), .B0(n1307), .B1(\rf<10><13> ), 
        .Y(n1523) );
  OAI221XL U484 ( .A0(n4154), .A1(n5162), .B0(n3994), .B1(n1304), .C0(n1515), 
        .Y(n1508) );
  AOI22X1 U485 ( .A0(n1306), .A1(\r15<14> ), .B0(n5155), .B1(\rf<10><14> ), 
        .Y(n1515) );
  OAI221XL U486 ( .A0(n4135), .A1(n5162), .B0(n3975), .B1(n1304), .C0(n1507), 
        .Y(n1500) );
  AOI22X1 U487 ( .A0(n1306), .A1(\r15<15> ), .B0(n5155), .B1(\rf<10><15> ), 
        .Y(n1507) );
  OAI221XL U488 ( .A0(n5195), .A1(n5267), .B0(n5192), .B1(n5093), .C0(n1255), 
        .Y(n1248) );
  AOI22X1 U489 ( .A0(n5191), .A1(n4645), .B0(n5188), .B1(n4869), .Y(n1255) );
  INVX1 U490 ( .A(\r15<12> ), .Y(n5267) );
  OAI221XL U491 ( .A0(n5195), .A1(n5266), .B0(n5192), .B1(n5094), .C0(n1247), 
        .Y(n1240) );
  AOI22X1 U492 ( .A0(n5190), .A1(n4646), .B0(n5188), .B1(n4870), .Y(n1247) );
  INVX1 U493 ( .A(\r15<13> ), .Y(n5266) );
  OAI221XL U494 ( .A0(n5195), .A1(n5265), .B0(n5192), .B1(n5095), .C0(n1239), 
        .Y(n1232) );
  AOI22X1 U495 ( .A0(n5191), .A1(n4647), .B0(n5188), .B1(n4871), .Y(n1239) );
  INVX1 U496 ( .A(\r15<14> ), .Y(n5265) );
  OAI221XL U497 ( .A0(n5195), .A1(n5264), .B0(n5192), .B1(n5096), .C0(n1231), 
        .Y(n1224) );
  AOI22X1 U498 ( .A0(n5190), .A1(n4648), .B0(n5188), .B1(n4872), .Y(n1231) );
  INVX1 U499 ( .A(\r15<15> ), .Y(n5264) );
  OAI221XL U500 ( .A0(n5195), .A1(n5263), .B0(n5192), .B1(n5097), .C0(n1223), 
        .Y(n1216) );
  AOI22X1 U501 ( .A0(n5191), .A1(n4649), .B0(n5188), .B1(n4873), .Y(n1223) );
  INVX1 U502 ( .A(\r15<16> ), .Y(n5263) );
  OR4X2 U503 ( .A(n1532), .B(n1533), .C(n1534), .D(n1535), .Y(\rd1<11> ) );
  OAI221XL U504 ( .A0(n4160), .A1(n5170), .B0(n4000), .B1(n5168), .C0(n1538), 
        .Y(n1533) );
  OAI221XL U505 ( .A0(n4161), .A1(n5178), .B0(n4001), .B1(n5176), .C0(n1537), 
        .Y(n1534) );
  OAI221XL U506 ( .A0(n4334), .A1(n5186), .B0(n4302), .B1(n5184), .C0(n1536), 
        .Y(n1535) );
  OR4X2 U507 ( .A(n1524), .B(n1525), .C(n1526), .D(n1527), .Y(\rd1<12> ) );
  OAI221XL U508 ( .A0(n4162), .A1(n5170), .B0(n4002), .B1(n5168), .C0(n1530), 
        .Y(n1525) );
  OAI221XL U509 ( .A0(n4163), .A1(n5178), .B0(n4003), .B1(n5176), .C0(n1529), 
        .Y(n1526) );
  OAI221XL U510 ( .A0(n4335), .A1(n5186), .B0(n4303), .B1(n5184), .C0(n1528), 
        .Y(n1527) );
  OR4X2 U511 ( .A(n1516), .B(n1517), .C(n1518), .D(n1519), .Y(\rd1<13> ) );
  OAI221XL U512 ( .A0(n4164), .A1(n5170), .B0(n4004), .B1(n5168), .C0(n1522), 
        .Y(n1517) );
  OAI221XL U513 ( .A0(n4165), .A1(n5178), .B0(n4005), .B1(n5176), .C0(n1521), 
        .Y(n1518) );
  OAI221XL U514 ( .A0(n4336), .A1(n5186), .B0(n4304), .B1(n5184), .C0(n1520), 
        .Y(n1519) );
  OR4X2 U515 ( .A(n1508), .B(n1509), .C(n1510), .D(n1511), .Y(\rd1<14> ) );
  OAI221XL U516 ( .A0(n4166), .A1(n5170), .B0(n4006), .B1(n5168), .C0(n1514), 
        .Y(n1509) );
  OAI221XL U517 ( .A0(n4167), .A1(n5178), .B0(n4007), .B1(n5176), .C0(n1513), 
        .Y(n1510) );
  OAI221XL U518 ( .A0(n4337), .A1(n5186), .B0(n4305), .B1(n5184), .C0(n1512), 
        .Y(n1511) );
  OR4X2 U519 ( .A(n1500), .B(n1501), .C(n1502), .D(n1503), .Y(\rd1<15> ) );
  OAI221XL U520 ( .A0(n4140), .A1(n5170), .B0(n3980), .B1(n5168), .C0(n1506), 
        .Y(n1501) );
  OAI221XL U521 ( .A0(n4141), .A1(n5178), .B0(n3981), .B1(n5176), .C0(n1505), 
        .Y(n1502) );
  OAI221XL U522 ( .A0(n4338), .A1(n5186), .B0(n4306), .B1(n5184), .C0(n1504), 
        .Y(n1503) );
  OAI221XL U523 ( .A0(n4150), .A1(n5162), .B0(n3990), .B1(n5159), .C0(n1547), 
        .Y(n1540) );
  AOI22X1 U524 ( .A0(n1306), .A1(\r15<10> ), .B0(n5155), .B1(\rf<10><10> ), 
        .Y(n1547) );
  OAI221XL U525 ( .A0(n5195), .A1(n5273), .B0(n5192), .B1(n5098), .C0(n1055), 
        .Y(n1048) );
  AOI22X1 U526 ( .A0(n5191), .A1(n4650), .B0(n5188), .B1(n4874), .Y(n1055) );
  INVX1 U527 ( .A(\r15<6> ), .Y(n5273) );
  OAI221XL U528 ( .A0(n5196), .A1(n5272), .B0(n5193), .B1(n5099), .C0(n1047), 
        .Y(n1040) );
  AOI22X1 U529 ( .A0(n5191), .A1(n4651), .B0(n5189), .B1(n4875), .Y(n1047) );
  INVX1 U530 ( .A(\r15<7> ), .Y(n5272) );
  OAI221XL U531 ( .A0(n5195), .A1(n5271), .B0(n5192), .B1(n5100), .C0(n1039), 
        .Y(n1032) );
  AOI22X1 U532 ( .A0(n5191), .A1(n4652), .B0(n5188), .B1(n4876), .Y(n1039) );
  INVX1 U533 ( .A(\r15<8> ), .Y(n5271) );
  OAI221XL U534 ( .A0(n5196), .A1(n5270), .B0(n5193), .B1(n5101), .C0(n1029), 
        .Y(n1008) );
  AOI22X1 U535 ( .A0(n5191), .A1(n4653), .B0(n5189), .B1(n4877), .Y(n1029) );
  INVX1 U536 ( .A(\r15<9> ), .Y(n5270) );
  OAI221XL U537 ( .A0(n5195), .A1(n5269), .B0(n5192), .B1(n5102), .C0(n1271), 
        .Y(n1264) );
  AOI22X1 U538 ( .A0(n5190), .A1(n4654), .B0(n5188), .B1(n4878), .Y(n1271) );
  INVX1 U539 ( .A(\r15<10> ), .Y(n5269) );
  OAI221XL U540 ( .A0(n5195), .A1(n5268), .B0(n5192), .B1(n5103), .C0(n1263), 
        .Y(n1256) );
  AOI22X1 U541 ( .A0(n5191), .A1(n4655), .B0(n5188), .B1(n4879), .Y(n1263) );
  INVX1 U542 ( .A(\r15<11> ), .Y(n5268) );
  OAI221XL U543 ( .A0(n4170), .A1(n5163), .B0(n4010), .B1(n5160), .C0(n1331), 
        .Y(n1324) );
  AOI22X1 U544 ( .A0(n1306), .A1(\r15<6> ), .B0(n1307), .B1(\rf<10><6> ), .Y(
        n1331) );
  OAI221XL U545 ( .A0(n4171), .A1(n5162), .B0(n4011), .B1(n5160), .C0(n1323), 
        .Y(n1316) );
  AOI22X1 U546 ( .A0(n1306), .A1(\r15<7> ), .B0(n1307), .B1(\rf<10><7> ), .Y(
        n1323) );
  OAI221XL U547 ( .A0(n4172), .A1(n5163), .B0(n4012), .B1(n5160), .C0(n1315), 
        .Y(n1308) );
  AOI22X1 U548 ( .A0(n1306), .A1(\r15<8> ), .B0(n1307), .B1(\rf<10><8> ), .Y(
        n1315) );
  OAI221XL U549 ( .A0(n4155), .A1(n5162), .B0(n3995), .B1(n5160), .C0(n1305), 
        .Y(n1284) );
  AOI22X1 U550 ( .A0(n1306), .A1(\r15<9> ), .B0(n1307), .B1(\rf<10><9> ), .Y(
        n1305) );
  OR4X2 U551 ( .A(n1324), .B(n1325), .C(n1326), .D(n1327), .Y(\rd1<6> ) );
  OAI221XL U552 ( .A0(n4177), .A1(n5171), .B0(n4017), .B1(n5169), .C0(n1330), 
        .Y(n1325) );
  OAI221XL U553 ( .A0(n4178), .A1(n5179), .B0(n4018), .B1(n5177), .C0(n1329), 
        .Y(n1326) );
  OAI221XL U554 ( .A0(n4329), .A1(n5187), .B0(n4297), .B1(n5185), .C0(n1328), 
        .Y(n1327) );
  OR4X2 U555 ( .A(n1316), .B(n1317), .C(n1318), .D(n1319), .Y(\rd1<7> ) );
  OAI221XL U556 ( .A0(n4179), .A1(n5170), .B0(n4019), .B1(n5168), .C0(n1322), 
        .Y(n1317) );
  OAI221XL U557 ( .A0(n4180), .A1(n5178), .B0(n4020), .B1(n5176), .C0(n1321), 
        .Y(n1318) );
  OAI221XL U558 ( .A0(n4330), .A1(n5186), .B0(n4298), .B1(n5184), .C0(n1320), 
        .Y(n1319) );
  OR4X2 U559 ( .A(n1308), .B(n1309), .C(n1310), .D(n1311), .Y(\rd1<8> ) );
  OAI221XL U560 ( .A0(n4181), .A1(n5171), .B0(n4021), .B1(n5169), .C0(n1314), 
        .Y(n1309) );
  OAI221XL U561 ( .A0(n4182), .A1(n5179), .B0(n4022), .B1(n5177), .C0(n1313), 
        .Y(n1310) );
  OAI221XL U562 ( .A0(n4331), .A1(n5187), .B0(n4299), .B1(n5185), .C0(n1312), 
        .Y(n1311) );
  OR4X2 U563 ( .A(n1284), .B(n1285), .C(n1286), .D(n1287), .Y(\rd1<9> ) );
  OAI221XL U564 ( .A0(n4156), .A1(n5170), .B0(n3996), .B1(n5168), .C0(n1300), 
        .Y(n1285) );
  OAI221XL U565 ( .A0(n4157), .A1(n5178), .B0(n3997), .B1(n5176), .C0(n1295), 
        .Y(n1286) );
  OAI221XL U566 ( .A0(n4332), .A1(n5186), .B0(n4300), .B1(n5184), .C0(n1290), 
        .Y(n1287) );
  OR4X2 U567 ( .A(n1540), .B(n1541), .C(n1542), .D(n1543), .Y(\rd1<10> ) );
  OAI221XL U568 ( .A0(n4158), .A1(n5170), .B0(n3998), .B1(n5168), .C0(n1546), 
        .Y(n1541) );
  OAI221XL U569 ( .A0(n4159), .A1(n5178), .B0(n3999), .B1(n5176), .C0(n1545), 
        .Y(n1542) );
  OAI221XL U570 ( .A0(n4333), .A1(n5186), .B0(n4301), .B1(n5184), .C0(n1544), 
        .Y(n1543) );
  OAI221XL U571 ( .A0(n4184), .A1(n5162), .B0(n4024), .B1(n5159), .C0(n1467), 
        .Y(n1460) );
  AOI22X1 U572 ( .A0(n1306), .A1(\r15<1> ), .B0(n5155), .B1(\rf<10><1> ), .Y(
        n1467) );
  OAI221XL U573 ( .A0(n4185), .A1(n5163), .B0(n4025), .B1(n5159), .C0(n1379), 
        .Y(n1372) );
  AOI22X1 U574 ( .A0(n5157), .A1(\r15<2> ), .B0(n5155), .B1(\rf<10><2> ), .Y(
        n1379) );
  OAI221XL U575 ( .A0(n4186), .A1(n5163), .B0(n4026), .B1(n5159), .C0(n1355), 
        .Y(n1348) );
  AOI22X1 U576 ( .A0(n5157), .A1(\r15<3> ), .B0(n1307), .B1(\rf<10><3> ), .Y(
        n1355) );
  OAI221XL U577 ( .A0(n5195), .A1(n5278), .B0(n5192), .B1(n5104), .C0(n1191), 
        .Y(n1184) );
  AOI22X1 U578 ( .A0(n5190), .A1(n4656), .B0(n5188), .B1(n4880), .Y(n1191) );
  INVX1 U579 ( .A(\r15<1> ), .Y(n5278) );
  OAI221XL U580 ( .A0(n5196), .A1(n5277), .B0(n5193), .B1(n5105), .C0(n1103), 
        .Y(n1096) );
  AOI22X1 U581 ( .A0(n5190), .A1(n4657), .B0(n5189), .B1(n4881), .Y(n1103) );
  INVX1 U582 ( .A(\r15<2> ), .Y(n5277) );
  OAI221XL U583 ( .A0(n5195), .A1(n5276), .B0(n5192), .B1(n5106), .C0(n1079), 
        .Y(n1072) );
  AOI22X1 U584 ( .A0(n5191), .A1(n4658), .B0(n5188), .B1(n4882), .Y(n1079) );
  INVX1 U585 ( .A(\r15<3> ), .Y(n5276) );
  OAI221XL U586 ( .A0(n5196), .A1(n5275), .B0(n1028), .B1(n5107), .C0(n1071), 
        .Y(n1064) );
  AOI22X1 U587 ( .A0(n5191), .A1(n4659), .B0(n5189), .B1(n4883), .Y(n1071) );
  INVX1 U588 ( .A(\r15<4> ), .Y(n5275) );
  OAI221XL U589 ( .A0(n5195), .A1(n5274), .B0(n1028), .B1(n5108), .C0(n1063), 
        .Y(n1056) );
  AOI22X1 U590 ( .A0(n5191), .A1(n4660), .B0(n5188), .B1(n4884), .Y(n1063) );
  INVX1 U591 ( .A(\r15<5> ), .Y(n5274) );
  OAI221XL U592 ( .A0(n4168), .A1(n5163), .B0(n4008), .B1(n5160), .C0(n1347), 
        .Y(n1340) );
  AOI22X1 U593 ( .A0(n5157), .A1(\r15<4> ), .B0(n1307), .B1(\rf<10><4> ), .Y(
        n1347) );
  OAI221XL U594 ( .A0(n4169), .A1(n5162), .B0(n4009), .B1(n5160), .C0(n1339), 
        .Y(n1332) );
  AOI22X1 U595 ( .A0(n5157), .A1(\r15<5> ), .B0(n1307), .B1(\rf<10><5> ), .Y(
        n1339) );
  OR4X2 U596 ( .A(n1460), .B(n1461), .C(n1462), .D(n1463), .Y(\rd1<1> ) );
  OAI221XL U597 ( .A0(n4189), .A1(n5170), .B0(n4029), .B1(n5168), .C0(n1466), 
        .Y(n1461) );
  OAI221XL U598 ( .A0(n4190), .A1(n5178), .B0(n4030), .B1(n5176), .C0(n1465), 
        .Y(n1462) );
  OAI221XL U599 ( .A0(n4324), .A1(n5186), .B0(n4292), .B1(n5184), .C0(n1464), 
        .Y(n1463) );
  OR4X2 U600 ( .A(n1372), .B(n1373), .C(n1374), .D(n1375), .Y(\rd1<2> ) );
  OAI221XL U601 ( .A0(n4191), .A1(n5171), .B0(n4031), .B1(n5169), .C0(n1378), 
        .Y(n1373) );
  OAI221XL U602 ( .A0(n4192), .A1(n5179), .B0(n4032), .B1(n5177), .C0(n1377), 
        .Y(n1374) );
  OAI221XL U603 ( .A0(n4325), .A1(n5187), .B0(n4293), .B1(n5185), .C0(n1376), 
        .Y(n1375) );
  OR4X2 U604 ( .A(n1348), .B(n1349), .C(n1350), .D(n1351), .Y(\rd1<3> ) );
  OAI221XL U605 ( .A0(n4193), .A1(n5171), .B0(n4033), .B1(n5169), .C0(n1354), 
        .Y(n1349) );
  OAI221XL U606 ( .A0(n4194), .A1(n5179), .B0(n4034), .B1(n5177), .C0(n1353), 
        .Y(n1350) );
  OAI221XL U607 ( .A0(n4326), .A1(n5187), .B0(n4294), .B1(n5185), .C0(n1352), 
        .Y(n1351) );
  OR4X2 U608 ( .A(n1340), .B(n1341), .C(n1342), .D(n1343), .Y(\rd1<4> ) );
  OAI221XL U609 ( .A0(n4173), .A1(n5171), .B0(n4013), .B1(n5169), .C0(n1346), 
        .Y(n1341) );
  OAI221XL U610 ( .A0(n4174), .A1(n5179), .B0(n4014), .B1(n5177), .C0(n1345), 
        .Y(n1342) );
  OAI221XL U611 ( .A0(n4327), .A1(n5187), .B0(n4295), .B1(n5185), .C0(n1344), 
        .Y(n1343) );
  OR4X2 U612 ( .A(n1332), .B(n1333), .C(n1334), .D(n1335), .Y(\rd1<5> ) );
  OAI221XL U613 ( .A0(n4175), .A1(n5170), .B0(n4015), .B1(n5168), .C0(n1338), 
        .Y(n1333) );
  OAI221XL U614 ( .A0(n4176), .A1(n5178), .B0(n4016), .B1(n5176), .C0(n1337), 
        .Y(n1334) );
  OAI221XL U615 ( .A0(n4328), .A1(n5186), .B0(n4296), .B1(n5184), .C0(n1336), 
        .Y(n1335) );
  OAI221XL U616 ( .A0(n4183), .A1(n5162), .B0(n4023), .B1(n5159), .C0(n1563), 
        .Y(n1548) );
  AOI22X1 U617 ( .A0(n1306), .A1(\r15<0> ), .B0(n5155), .B1(\rf<10><0> ), .Y(
        n1563) );
  OAI221XL U618 ( .A0(n5195), .A1(n5279), .B0(n5192), .B1(n5109), .C0(n1283), 
        .Y(n1272) );
  AOI22X1 U619 ( .A0(n5191), .A1(n4661), .B0(n5188), .B1(n4885), .Y(n1283) );
  INVX1 U620 ( .A(\r15<0> ), .Y(n5279) );
  OR4X2 U621 ( .A(n1548), .B(n1549), .C(n1550), .D(n1551), .Y(\rd1<0> ) );
  OAI221XL U622 ( .A0(n4187), .A1(n5170), .B0(n4027), .B1(n5168), .C0(n1561), 
        .Y(n1549) );
  OAI221XL U623 ( .A0(n4188), .A1(n5178), .B0(n4028), .B1(n5176), .C0(n1559), 
        .Y(n1550) );
  OAI221XL U624 ( .A0(n4323), .A1(n5186), .B0(n4291), .B1(n5184), .C0(n1552), 
        .Y(n1551) );
  NAND3X1 U625 ( .A(we3), .B(n5287), .C(\wa3<3> ), .Y(n1568) );
  NAND3X1 U626 ( .A(we3), .B(n5285), .C(\wa3<0> ), .Y(n1570) );
  NAND3X1 U627 ( .A(\wa3<3> ), .B(we3), .C(\wa3<0> ), .Y(n1569) );
  AOI22X1 U628 ( .A0(n5182), .A1(n4387), .B0(n5180), .B1(n4355), .Y(n1552) );
  AOI22X1 U629 ( .A0(n5174), .A1(\rf<7><0> ), .B0(n1297), .B1(\rf<2><0> ), .Y(
        n1559) );
  AOI22X1 U630 ( .A0(n5166), .A1(\rf<11><0> ), .B0(n5164), .B1(\rf<6><0> ), 
        .Y(n1561) );
  AOI22X1 U631 ( .A0(n1291), .A1(n4388), .B0(n5180), .B1(n4356), .Y(n1464) );
  AOI22X1 U632 ( .A0(n5174), .A1(\rf<7><1> ), .B0(n1297), .B1(\rf<2><1> ), .Y(
        n1465) );
  AOI22X1 U633 ( .A0(n5166), .A1(\rf<11><1> ), .B0(n5164), .B1(\rf<6><1> ), 
        .Y(n1466) );
  AOI22X1 U634 ( .A0(n5182), .A1(n4389), .B0(n1292), .B1(n4357), .Y(n1376) );
  AOI22X1 U635 ( .A0(n1296), .A1(\rf<7><2> ), .B0(n5172), .B1(\rf<2><2> ), .Y(
        n1377) );
  AOI22X1 U636 ( .A0(n5166), .A1(\rf<11><2> ), .B0(n1302), .B1(\rf<6><2> ), 
        .Y(n1378) );
  AOI22X1 U637 ( .A0(n1291), .A1(n4390), .B0(n1292), .B1(n4358), .Y(n1352) );
  AOI22X1 U638 ( .A0(n1296), .A1(\rf<7><3> ), .B0(n1297), .B1(\rf<2><3> ), .Y(
        n1353) );
  AOI22X1 U639 ( .A0(n5166), .A1(\rf<11><3> ), .B0(n1302), .B1(\rf<6><3> ), 
        .Y(n1354) );
  AOI22X1 U640 ( .A0(n1291), .A1(n4391), .B0(n1292), .B1(n4359), .Y(n1344) );
  AOI22X1 U641 ( .A0(n1296), .A1(\rf<7><4> ), .B0(n5172), .B1(\rf<2><4> ), .Y(
        n1345) );
  AOI22X1 U642 ( .A0(n1301), .A1(\rf<11><4> ), .B0(n1302), .B1(\rf<6><4> ), 
        .Y(n1346) );
  AOI22X1 U643 ( .A0(n1291), .A1(n4392), .B0(n1292), .B1(n4360), .Y(n1336) );
  AOI22X1 U644 ( .A0(n1296), .A1(\rf<7><5> ), .B0(n5172), .B1(\rf<2><5> ), .Y(
        n1337) );
  AOI22X1 U645 ( .A0(n1301), .A1(\rf<11><5> ), .B0(n1302), .B1(\rf<6><5> ), 
        .Y(n1338) );
  AOI22X1 U646 ( .A0(n1291), .A1(n4393), .B0(n1292), .B1(n4361), .Y(n1328) );
  AOI22X1 U647 ( .A0(n1296), .A1(\rf<7><6> ), .B0(n1297), .B1(\rf<2><6> ), .Y(
        n1329) );
  AOI22X1 U648 ( .A0(n1301), .A1(\rf<11><6> ), .B0(n1302), .B1(\rf<6><6> ), 
        .Y(n1330) );
  AOI22X1 U649 ( .A0(n1291), .A1(n4394), .B0(n1292), .B1(n4362), .Y(n1320) );
  AOI22X1 U650 ( .A0(n1296), .A1(\rf<7><7> ), .B0(n1297), .B1(\rf<2><7> ), .Y(
        n1321) );
  AOI22X1 U651 ( .A0(n1301), .A1(\rf<11><7> ), .B0(n1302), .B1(\rf<6><7> ), 
        .Y(n1322) );
  AOI22X1 U652 ( .A0(n1291), .A1(n4395), .B0(n1292), .B1(n4363), .Y(n1312) );
  AOI22X1 U653 ( .A0(n1296), .A1(\rf<7><8> ), .B0(n1297), .B1(\rf<2><8> ), .Y(
        n1313) );
  AOI22X1 U654 ( .A0(n5166), .A1(\rf<11><8> ), .B0(n1302), .B1(\rf<6><8> ), 
        .Y(n1314) );
  AOI22X1 U655 ( .A0(n1291), .A1(n4396), .B0(n1292), .B1(n4364), .Y(n1290) );
  AOI22X1 U656 ( .A0(n1296), .A1(\rf<7><9> ), .B0(n1297), .B1(\rf<2><9> ), .Y(
        n1295) );
  AOI22X1 U657 ( .A0(n5166), .A1(\rf<11><9> ), .B0(n1302), .B1(\rf<6><9> ), 
        .Y(n1300) );
  AOI22X1 U658 ( .A0(n1291), .A1(n4397), .B0(n5180), .B1(n4365), .Y(n1544) );
  AOI22X1 U659 ( .A0(n5174), .A1(\rf<7><10> ), .B0(n1297), .B1(\rf<2><10> ), 
        .Y(n1545) );
  AOI22X1 U660 ( .A0(n5166), .A1(\rf<11><10> ), .B0(n5164), .B1(\rf<6><10> ), 
        .Y(n1546) );
  AOI22X1 U661 ( .A0(n1291), .A1(n4398), .B0(n5180), .B1(n4366), .Y(n1536) );
  AOI22X1 U662 ( .A0(n5174), .A1(\rf<7><11> ), .B0(n1297), .B1(\rf<2><11> ), 
        .Y(n1537) );
  AOI22X1 U663 ( .A0(n5166), .A1(\rf<11><11> ), .B0(n5164), .B1(\rf<6><11> ), 
        .Y(n1538) );
  AOI22X1 U664 ( .A0(n1291), .A1(n4399), .B0(n5180), .B1(n4367), .Y(n1528) );
  AOI22X1 U665 ( .A0(n5174), .A1(\rf<7><12> ), .B0(n1297), .B1(\rf<2><12> ), 
        .Y(n1529) );
  AOI22X1 U666 ( .A0(n1301), .A1(\rf<11><12> ), .B0(n5164), .B1(\rf<6><12> ), 
        .Y(n1530) );
  AOI22X1 U667 ( .A0(n5182), .A1(n4400), .B0(n5180), .B1(n4368), .Y(n1520) );
  AOI22X1 U668 ( .A0(n5174), .A1(\rf<7><13> ), .B0(n1297), .B1(\rf<2><13> ), 
        .Y(n1521) );
  AOI22X1 U669 ( .A0(n1301), .A1(\rf<11><13> ), .B0(n5164), .B1(\rf<6><13> ), 
        .Y(n1522) );
  AOI22X1 U670 ( .A0(n5182), .A1(n4401), .B0(n5180), .B1(n4369), .Y(n1512) );
  AOI22X1 U671 ( .A0(n5174), .A1(\rf<7><14> ), .B0(n1297), .B1(\rf<2><14> ), 
        .Y(n1513) );
  AOI22X1 U672 ( .A0(n1301), .A1(\rf<11><14> ), .B0(n5164), .B1(\rf<6><14> ), 
        .Y(n1514) );
  AOI22X1 U673 ( .A0(n5182), .A1(n4402), .B0(n5180), .B1(n4370), .Y(n1504) );
  AOI22X1 U674 ( .A0(n5174), .A1(\rf<7><15> ), .B0(n5172), .B1(\rf<2><15> ), 
        .Y(n1505) );
  AOI22X1 U675 ( .A0(n1301), .A1(\rf<11><15> ), .B0(n5164), .B1(\rf<6><15> ), 
        .Y(n1506) );
  AOI22X1 U676 ( .A0(n5182), .A1(n4403), .B0(n5180), .B1(n4371), .Y(n1496) );
  AOI22X1 U677 ( .A0(n5174), .A1(\rf<7><16> ), .B0(n5172), .B1(\rf<2><16> ), 
        .Y(n1497) );
  AOI22X1 U678 ( .A0(n1301), .A1(\rf<11><16> ), .B0(n5164), .B1(\rf<6><16> ), 
        .Y(n1498) );
  AOI22X1 U679 ( .A0(n5182), .A1(n4404), .B0(n5180), .B1(n4372), .Y(n1488) );
  AOI22X1 U680 ( .A0(n5174), .A1(\rf<7><17> ), .B0(n5172), .B1(\rf<2><17> ), 
        .Y(n1489) );
  AOI22X1 U681 ( .A0(n1301), .A1(\rf<11><17> ), .B0(n5164), .B1(\rf<6><17> ), 
        .Y(n1490) );
  AOI22X1 U682 ( .A0(n5182), .A1(n4405), .B0(n5180), .B1(n4373), .Y(n1480) );
  AOI22X1 U683 ( .A0(n5174), .A1(\rf<7><18> ), .B0(n5172), .B1(\rf<2><18> ), 
        .Y(n1481) );
  AOI22X1 U684 ( .A0(n1301), .A1(\rf<11><18> ), .B0(n5164), .B1(\rf<6><18> ), 
        .Y(n1482) );
  AOI22X1 U685 ( .A0(n5182), .A1(n4406), .B0(n5180), .B1(n4374), .Y(n1472) );
  AOI22X1 U686 ( .A0(n5174), .A1(\rf<7><19> ), .B0(n5172), .B1(\rf<2><19> ), 
        .Y(n1473) );
  AOI22X1 U687 ( .A0(n1301), .A1(\rf<11><19> ), .B0(n5164), .B1(\rf<6><19> ), 
        .Y(n1474) );
  AOI22X1 U688 ( .A0(n5182), .A1(n4407), .B0(n1292), .B1(n4375), .Y(n1456) );
  AOI22X1 U689 ( .A0(n1296), .A1(\rf<7><20> ), .B0(n5172), .B1(\rf<2><20> ), 
        .Y(n1457) );
  AOI22X1 U690 ( .A0(n5166), .A1(\rf<11><20> ), .B0(n1302), .B1(\rf<6><20> ), 
        .Y(n1458) );
  AOI22X1 U691 ( .A0(n5182), .A1(n4408), .B0(n1292), .B1(n4376), .Y(n1448) );
  AOI22X1 U692 ( .A0(n1296), .A1(\rf<7><21> ), .B0(n5172), .B1(\rf<2><21> ), 
        .Y(n1449) );
  AOI22X1 U693 ( .A0(n5166), .A1(\rf<11><21> ), .B0(n1302), .B1(\rf<6><21> ), 
        .Y(n1450) );
  AOI22X1 U694 ( .A0(n5182), .A1(n4409), .B0(n1292), .B1(n4377), .Y(n1440) );
  AOI22X1 U695 ( .A0(n1296), .A1(\rf<7><22> ), .B0(n5172), .B1(\rf<2><22> ), 
        .Y(n1441) );
  AOI22X1 U696 ( .A0(n5166), .A1(\rf<11><22> ), .B0(n1302), .B1(\rf<6><22> ), 
        .Y(n1442) );
  AOI22X1 U697 ( .A0(n5182), .A1(n4410), .B0(n1292), .B1(n4378), .Y(n1432) );
  AOI22X1 U698 ( .A0(n5174), .A1(\rf<7><23> ), .B0(n5172), .B1(\rf<2><23> ), 
        .Y(n1433) );
  AOI22X1 U699 ( .A0(n5166), .A1(\rf<11><23> ), .B0(n1302), .B1(\rf<6><23> ), 
        .Y(n1434) );
  AOI22X1 U700 ( .A0(n5182), .A1(n4411), .B0(n5180), .B1(n4379), .Y(n1424) );
  AOI22X1 U701 ( .A0(n5174), .A1(\rf<7><24> ), .B0(n5172), .B1(\rf<2><24> ), 
        .Y(n1425) );
  AOI22X1 U702 ( .A0(n5166), .A1(\rf<11><24> ), .B0(n5164), .B1(\rf<6><24> ), 
        .Y(n1426) );
  AOI22X1 U703 ( .A0(n5182), .A1(n4412), .B0(n5180), .B1(n4380), .Y(n1416) );
  AOI22X1 U704 ( .A0(n5174), .A1(\rf<7><25> ), .B0(n5172), .B1(\rf<2><25> ), 
        .Y(n1417) );
  AOI22X1 U705 ( .A0(n5166), .A1(\rf<11><25> ), .B0(n5164), .B1(\rf<6><25> ), 
        .Y(n1418) );
  AOI22X1 U706 ( .A0(n5182), .A1(n4413), .B0(n5180), .B1(n4381), .Y(n1408) );
  AOI22X1 U707 ( .A0(n5174), .A1(\rf<7><26> ), .B0(n5172), .B1(\rf<2><26> ), 
        .Y(n1409) );
  AOI22X1 U708 ( .A0(n5166), .A1(\rf<11><26> ), .B0(n5164), .B1(\rf<6><26> ), 
        .Y(n1410) );
  AOI22X1 U709 ( .A0(n5182), .A1(n4414), .B0(n5180), .B1(n4382), .Y(n1400) );
  AOI22X1 U710 ( .A0(n5174), .A1(\rf<7><27> ), .B0(n5172), .B1(\rf<2><27> ), 
        .Y(n1401) );
  AOI22X1 U711 ( .A0(n5166), .A1(\rf<11><27> ), .B0(n5164), .B1(\rf<6><27> ), 
        .Y(n1402) );
  AOI22X1 U712 ( .A0(n5182), .A1(n4415), .B0(n5180), .B1(n4383), .Y(n1392) );
  AOI22X1 U713 ( .A0(n5174), .A1(\rf<7><28> ), .B0(n5172), .B1(\rf<2><28> ), 
        .Y(n1393) );
  AOI22X1 U714 ( .A0(n5166), .A1(\rf<11><28> ), .B0(n5164), .B1(\rf<6><28> ), 
        .Y(n1394) );
  AOI22X1 U715 ( .A0(n5182), .A1(n4416), .B0(n5180), .B1(n4384), .Y(n1384) );
  AOI22X1 U716 ( .A0(n5174), .A1(\rf<7><29> ), .B0(n5172), .B1(\rf<2><29> ), 
        .Y(n1385) );
  AOI22X1 U717 ( .A0(n5166), .A1(\rf<11><29> ), .B0(n5164), .B1(\rf<6><29> ), 
        .Y(n1386) );
  AOI22X1 U718 ( .A0(n5182), .A1(n4417), .B0(n5180), .B1(n4385), .Y(n1368) );
  AOI22X1 U719 ( .A0(n5174), .A1(\rf<7><30> ), .B0(n5172), .B1(\rf<2><30> ), 
        .Y(n1369) );
  AOI22X1 U720 ( .A0(n5166), .A1(\rf<11><30> ), .B0(n5164), .B1(\rf<6><30> ), 
        .Y(n1370) );
  AOI22X1 U721 ( .A0(n1291), .A1(n4418), .B0(n1292), .B1(n4386), .Y(n1360) );
  AOI22X1 U722 ( .A0(n1296), .A1(\rf<7><31> ), .B0(n1297), .B1(\rf<2><31> ), 
        .Y(n1361) );
  AOI22X1 U723 ( .A0(n5166), .A1(\rf<11><31> ), .B0(n1302), .B1(\rf<6><31> ), 
        .Y(n1362) );
  AOI22X1 U724 ( .A0(n5215), .A1(n4662), .B0(n5213), .B1(n4886), .Y(n1276) );
  AOI22X1 U725 ( .A0(n5199), .A1(n4663), .B0(n5197), .B1(n4887), .Y(n1282) );
  AOI22X1 U726 ( .A0(n5207), .A1(n4664), .B0(n5205), .B1(n4888), .Y(n1280) );
  AOI22X1 U727 ( .A0(n5215), .A1(n4665), .B0(n5213), .B1(n4889), .Y(n1188) );
  AOI22X1 U728 ( .A0(n5199), .A1(n4666), .B0(n5197), .B1(n4890), .Y(n1190) );
  AOI22X1 U729 ( .A0(n5207), .A1(n4667), .B0(n5205), .B1(n4891), .Y(n1189) );
  AOI22X1 U730 ( .A0(n5216), .A1(n4668), .B0(n5214), .B1(n4892), .Y(n1100) );
  AOI22X1 U731 ( .A0(n5200), .A1(n4669), .B0(n5198), .B1(n4893), .Y(n1102) );
  AOI22X1 U732 ( .A0(n5208), .A1(n4670), .B0(n5206), .B1(n4894), .Y(n1101) );
  AOI22X1 U733 ( .A0(n5216), .A1(n4671), .B0(n5214), .B1(n4895), .Y(n1076) );
  AOI22X1 U734 ( .A0(n5200), .A1(n4672), .B0(n5198), .B1(n4896), .Y(n1078) );
  AOI22X1 U735 ( .A0(n5208), .A1(n4673), .B0(n5206), .B1(n4897), .Y(n1077) );
  AOI22X1 U736 ( .A0(n5216), .A1(n4674), .B0(n5213), .B1(n4898), .Y(n1068) );
  AOI22X1 U737 ( .A0(n5200), .A1(n4675), .B0(n5197), .B1(n4899), .Y(n1070) );
  AOI22X1 U738 ( .A0(n5208), .A1(n4676), .B0(n5205), .B1(n4900), .Y(n1069) );
  AOI22X1 U739 ( .A0(n5216), .A1(n4677), .B0(n5214), .B1(n4901), .Y(n1060) );
  AOI22X1 U740 ( .A0(n5200), .A1(n4678), .B0(n5198), .B1(n4902), .Y(n1062) );
  AOI22X1 U741 ( .A0(n5208), .A1(n4679), .B0(n5206), .B1(n4903), .Y(n1061) );
  AOI22X1 U742 ( .A0(n5216), .A1(n4680), .B0(n5213), .B1(n4904), .Y(n1052) );
  AOI22X1 U743 ( .A0(n5200), .A1(n4681), .B0(n5197), .B1(n4905), .Y(n1054) );
  AOI22X1 U744 ( .A0(n5208), .A1(n4682), .B0(n5205), .B1(n4906), .Y(n1053) );
  AOI22X1 U745 ( .A0(n5216), .A1(n4683), .B0(n5214), .B1(n4907), .Y(n1044) );
  AOI22X1 U746 ( .A0(n5200), .A1(n4684), .B0(n5198), .B1(n4908), .Y(n1046) );
  AOI22X1 U747 ( .A0(n5208), .A1(n4685), .B0(n5206), .B1(n4909), .Y(n1045) );
  AOI22X1 U748 ( .A0(n5216), .A1(n4686), .B0(n5213), .B1(n4910), .Y(n1036) );
  AOI22X1 U749 ( .A0(n5200), .A1(n4687), .B0(n5197), .B1(n4911), .Y(n1038) );
  AOI22X1 U750 ( .A0(n5208), .A1(n4688), .B0(n5205), .B1(n4912), .Y(n1037) );
  AOI22X1 U751 ( .A0(n5216), .A1(n4689), .B0(n5214), .B1(n4913), .Y(n1014) );
  AOI22X1 U752 ( .A0(n5200), .A1(n4690), .B0(n5198), .B1(n4914), .Y(n1024) );
  AOI22X1 U753 ( .A0(n5208), .A1(n4691), .B0(n5206), .B1(n4915), .Y(n1019) );
  AOI22X1 U754 ( .A0(n5215), .A1(n4692), .B0(n5213), .B1(n4916), .Y(n1268) );
  AOI22X1 U755 ( .A0(n5199), .A1(n4693), .B0(n5197), .B1(n4917), .Y(n1270) );
  AOI22X1 U756 ( .A0(n5207), .A1(n4694), .B0(n5205), .B1(n4918), .Y(n1269) );
  AOI22X1 U757 ( .A0(n5215), .A1(n4695), .B0(n5213), .B1(n4919), .Y(n1260) );
  AOI22X1 U758 ( .A0(n5199), .A1(n4696), .B0(n5197), .B1(n4920), .Y(n1262) );
  AOI22X1 U759 ( .A0(n5207), .A1(n4697), .B0(n5205), .B1(n4921), .Y(n1261) );
  AOI22X1 U760 ( .A0(n5215), .A1(n4698), .B0(n5213), .B1(n4922), .Y(n1252) );
  AOI22X1 U761 ( .A0(n5199), .A1(n4699), .B0(n5197), .B1(n4923), .Y(n1254) );
  AOI22X1 U762 ( .A0(n5207), .A1(n4700), .B0(n5205), .B1(n4924), .Y(n1253) );
  AOI22X1 U763 ( .A0(n5215), .A1(n4701), .B0(n5213), .B1(n4925), .Y(n1244) );
  AOI22X1 U764 ( .A0(n5199), .A1(n4702), .B0(n5197), .B1(n4926), .Y(n1246) );
  AOI22X1 U765 ( .A0(n5207), .A1(n4703), .B0(n5205), .B1(n4927), .Y(n1245) );
  AOI22X1 U766 ( .A0(n5215), .A1(n4704), .B0(n5213), .B1(n4928), .Y(n1236) );
  AOI22X1 U767 ( .A0(n5199), .A1(n4705), .B0(n5197), .B1(n4929), .Y(n1238) );
  AOI22X1 U768 ( .A0(n5207), .A1(n4706), .B0(n5205), .B1(n4930), .Y(n1237) );
  AOI22X1 U769 ( .A0(n5215), .A1(n4707), .B0(n5213), .B1(n4931), .Y(n1228) );
  AOI22X1 U770 ( .A0(n5199), .A1(n4708), .B0(n5197), .B1(n4932), .Y(n1230) );
  AOI22X1 U771 ( .A0(n5207), .A1(n4709), .B0(n5205), .B1(n4933), .Y(n1229) );
  AOI22X1 U772 ( .A0(n5215), .A1(n4710), .B0(n5213), .B1(n4934), .Y(n1220) );
  AOI22X1 U773 ( .A0(n5199), .A1(n4711), .B0(n5197), .B1(n4935), .Y(n1222) );
  AOI22X1 U774 ( .A0(n5207), .A1(n4712), .B0(n5205), .B1(n4936), .Y(n1221) );
  AOI22X1 U775 ( .A0(n5215), .A1(n4713), .B0(n5213), .B1(n4937), .Y(n1212) );
  AOI22X1 U776 ( .A0(n5199), .A1(n4714), .B0(n5197), .B1(n4938), .Y(n1214) );
  AOI22X1 U777 ( .A0(n5207), .A1(n4715), .B0(n5205), .B1(n4939), .Y(n1213) );
  AOI22X1 U778 ( .A0(n5215), .A1(n4716), .B0(n5213), .B1(n4940), .Y(n1204) );
  AOI22X1 U779 ( .A0(n5199), .A1(n4717), .B0(n5197), .B1(n4941), .Y(n1206) );
  AOI22X1 U780 ( .A0(n5207), .A1(n4718), .B0(n5205), .B1(n4942), .Y(n1205) );
  AOI22X1 U781 ( .A0(n5215), .A1(n4719), .B0(n5213), .B1(n4943), .Y(n1196) );
  AOI22X1 U782 ( .A0(n5199), .A1(n4720), .B0(n5197), .B1(n4944), .Y(n1198) );
  AOI22X1 U783 ( .A0(n5207), .A1(n4721), .B0(n5205), .B1(n4945), .Y(n1197) );
  AOI22X1 U784 ( .A0(n5216), .A1(n4722), .B0(n5214), .B1(n4946), .Y(n1180) );
  AOI22X1 U785 ( .A0(n5200), .A1(n4723), .B0(n5198), .B1(n4947), .Y(n1182) );
  AOI22X1 U786 ( .A0(n5208), .A1(n4724), .B0(n5206), .B1(n4948), .Y(n1181) );
  AOI22X1 U787 ( .A0(n5216), .A1(n4725), .B0(n5214), .B1(n4949), .Y(n1172) );
  AOI22X1 U788 ( .A0(n5200), .A1(n4726), .B0(n5198), .B1(n4950), .Y(n1174) );
  AOI22X1 U789 ( .A0(n5208), .A1(n4727), .B0(n5206), .B1(n4951), .Y(n1173) );
  AOI22X1 U790 ( .A0(n5216), .A1(n4728), .B0(n5214), .B1(n4952), .Y(n1164) );
  AOI22X1 U791 ( .A0(n5200), .A1(n4729), .B0(n5198), .B1(n4953), .Y(n1166) );
  AOI22X1 U792 ( .A0(n5208), .A1(n4730), .B0(n5206), .B1(n4954), .Y(n1165) );
  AOI22X1 U793 ( .A0(n5215), .A1(n4731), .B0(n5214), .B1(n4955), .Y(n1156) );
  AOI22X1 U794 ( .A0(n5199), .A1(n4732), .B0(n5198), .B1(n4956), .Y(n1158) );
  AOI22X1 U795 ( .A0(n5207), .A1(n4733), .B0(n5206), .B1(n4957), .Y(n1157) );
  AOI22X1 U796 ( .A0(n5216), .A1(n4734), .B0(n5214), .B1(n4958), .Y(n1148) );
  AOI22X1 U797 ( .A0(n5200), .A1(n4735), .B0(n5198), .B1(n4959), .Y(n1150) );
  AOI22X1 U798 ( .A0(n5208), .A1(n4736), .B0(n5206), .B1(n4960), .Y(n1149) );
  AOI22X1 U799 ( .A0(n5215), .A1(n4737), .B0(n5214), .B1(n4961), .Y(n1140) );
  AOI22X1 U800 ( .A0(n5199), .A1(n4738), .B0(n5198), .B1(n4962), .Y(n1142) );
  AOI22X1 U801 ( .A0(n5207), .A1(n4739), .B0(n5206), .B1(n4963), .Y(n1141) );
  AOI22X1 U802 ( .A0(n5216), .A1(n4740), .B0(n5214), .B1(n4964), .Y(n1132) );
  AOI22X1 U803 ( .A0(n5200), .A1(n4741), .B0(n5198), .B1(n4965), .Y(n1134) );
  AOI22X1 U804 ( .A0(n5208), .A1(n4742), .B0(n5206), .B1(n4966), .Y(n1133) );
  AOI22X1 U805 ( .A0(n5215), .A1(n4743), .B0(n5214), .B1(n4967), .Y(n1124) );
  AOI22X1 U806 ( .A0(n5199), .A1(n4744), .B0(n5198), .B1(n4968), .Y(n1126) );
  AOI22X1 U807 ( .A0(n5207), .A1(n4745), .B0(n5206), .B1(n4969), .Y(n1125) );
  AOI22X1 U808 ( .A0(n5216), .A1(n4746), .B0(n5214), .B1(n4970), .Y(n1116) );
  AOI22X1 U809 ( .A0(n5200), .A1(n4747), .B0(n5198), .B1(n4971), .Y(n1118) );
  AOI22X1 U810 ( .A0(n5208), .A1(n4748), .B0(n5206), .B1(n4972), .Y(n1117) );
  AOI22X1 U811 ( .A0(n5215), .A1(n4749), .B0(n5214), .B1(n4973), .Y(n1108) );
  AOI22X1 U812 ( .A0(n5199), .A1(n4750), .B0(n5198), .B1(n4974), .Y(n1110) );
  AOI22X1 U813 ( .A0(n5207), .A1(n4751), .B0(n5206), .B1(n4975), .Y(n1109) );
  AOI22X1 U814 ( .A0(n5216), .A1(n4752), .B0(n5214), .B1(n4976), .Y(n1092) );
  AOI22X1 U815 ( .A0(n5200), .A1(n4753), .B0(n5198), .B1(n4977), .Y(n1094) );
  AOI22X1 U816 ( .A0(n5208), .A1(n4754), .B0(n5206), .B1(n4978), .Y(n1093) );
  AOI22X1 U817 ( .A0(n5216), .A1(n4755), .B0(n5213), .B1(n4979), .Y(n1084) );
  AOI22X1 U818 ( .A0(n5200), .A1(n4756), .B0(n5197), .B1(n4980), .Y(n1086) );
  AOI22X1 U819 ( .A0(n5208), .A1(n4757), .B0(n5205), .B1(n4981), .Y(n1085) );
  BUFX3 U820 ( .A(N16), .Y(n5142) );
  NAND2X1 U821 ( .A(\wa3<2> ), .B(n5289), .Y(n1567) );
  NAND2X1 U822 ( .A(\wa3<1> ), .B(n5283), .Y(n1565) );
  NAND2X1 U823 ( .A(\wa3<2> ), .B(\wa3<1> ), .Y(n1571) );
  INVX1 U824 ( .A(\wa3<1> ), .Y(n5289) );
  INVX1 U825 ( .A(\wa3<2> ), .Y(n5283) );
  INVX1 U826 ( .A(\wa3<3> ), .Y(n5285) );
  INVX1 U827 ( .A(\wa3<0> ), .Y(n5287) );
endmodule


module extend ( .Instr({\Instr<23> , \Instr<22> , \Instr<21> , \Instr<20> , 
        \Instr<19> , \Instr<18> , \Instr<17> , \Instr<16> , \Instr<15> , 
        \Instr<14> , \Instr<13> , \Instr<12> , \Instr<11> , \Instr<10> , 
        \Instr<9> , \Instr<8> , \Instr<7> , \Instr<6> , \Instr<5> , \Instr<4> , 
        \Instr<3> , \Instr<2> , \Instr<1> , \Instr<0> }), .ImmSrc({\ImmSrc<1> , 
        \ImmSrc<0> }), .ExtImm({\ExtImm<31> , \ExtImm<30> , \ExtImm<29> , 
        \ExtImm<28> , \ExtImm<27> , \ExtImm<26> , \ExtImm<25> , \ExtImm<24> , 
        \ExtImm<23> , \ExtImm<22> , \ExtImm<21> , \ExtImm<20> , \ExtImm<19> , 
        \ExtImm<18> , \ExtImm<17> , \ExtImm<16> , \ExtImm<15> , \ExtImm<14> , 
        \ExtImm<13> , \ExtImm<12> , \ExtImm<11> , \ExtImm<10> , \ExtImm<9> , 
        \ExtImm<8> , \ExtImm<7> , \ExtImm<6> , \ExtImm<5> , \ExtImm<4> , 
        \ExtImm<3> , \ExtImm<2> , \ExtImm<1> , \ExtImm<0> }) );
  input \Instr<23> , \Instr<22> , \Instr<21> , \Instr<20> , \Instr<19> ,
         \Instr<18> , \Instr<17> , \Instr<16> , \Instr<15> , \Instr<14> ,
         \Instr<13> , \Instr<12> , \Instr<11> , \Instr<10> , \Instr<9> ,
         \Instr<8> , \Instr<7> , \Instr<6> , \Instr<5> , \Instr<4> ,
         \Instr<3> , \Instr<2> , \Instr<1> , \Instr<0> , \ImmSrc<1> ,
         \ImmSrc<0> ;
  output \ExtImm<31> , \ExtImm<30> , \ExtImm<29> , \ExtImm<28> , \ExtImm<27> ,
         \ExtImm<26> , \ExtImm<25> , \ExtImm<24> , \ExtImm<23> , \ExtImm<22> ,
         \ExtImm<21> , \ExtImm<20> , \ExtImm<19> , \ExtImm<18> , \ExtImm<17> ,
         \ExtImm<16> , \ExtImm<15> , \ExtImm<14> , \ExtImm<13> , \ExtImm<12> ,
         \ExtImm<11> , \ExtImm<10> , \ExtImm<9> , \ExtImm<8> , \ExtImm<7> ,
         \ExtImm<6> , \ExtImm<5> , \ExtImm<4> , \ExtImm<3> , \ExtImm<2> ,
         \ExtImm<1> , \ExtImm<0> ;
  wire   n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151,
         n152, n153, n154, n155;

  BUFX3 U2 ( .A(n155), .Y(n141) );
  INVX1 U3 ( .A(\ImmSrc<1> ), .Y(n155) );
  NOR2X1 U4 ( .A(\ImmSrc<1> ), .B(n152), .Y(\ExtImm<1> ) );
  NOR2X1 U5 ( .A(\ImmSrc<1> ), .B(n153), .Y(\ExtImm<0> ) );
  OAI22X1 U6 ( .A0(n141), .A1(n153), .B0(\ImmSrc<1> ), .B1(n151), .Y(
        \ExtImm<2> ) );
  OAI22X1 U7 ( .A0(n141), .A1(n152), .B0(\ImmSrc<1> ), .B1(n150), .Y(
        \ExtImm<3> ) );
  OAI22X1 U8 ( .A0(n141), .A1(n151), .B0(\ImmSrc<1> ), .B1(n149), .Y(
        \ExtImm<4> ) );
  OAI22X1 U9 ( .A0(n141), .A1(n150), .B0(\ImmSrc<1> ), .B1(n148), .Y(
        \ExtImm<5> ) );
  OAI22X1 U10 ( .A0(n141), .A1(n149), .B0(\ImmSrc<1> ), .B1(n147), .Y(
        \ExtImm<6> ) );
  OAI22X1 U11 ( .A0(n141), .A1(n147), .B0(n154), .B1(n145), .Y(\ExtImm<8> ) );
  OAI22X1 U12 ( .A0(n141), .A1(n145), .B0(n154), .B1(n143), .Y(\ExtImm<10> )
         );
  OAI22X1 U13 ( .A0(n144), .A1(n141), .B0(n154), .B1(n142), .Y(\ExtImm<11> )
         );
  OAI22X1 U14 ( .A0(n141), .A1(n146), .B0(n154), .B1(n144), .Y(\ExtImm<9> ) );
  OAI22X1 U15 ( .A0(n141), .A1(n148), .B0(\ImmSrc<1> ), .B1(n146), .Y(
        \ExtImm<7> ) );
  NOR2BX1 U16 ( .AN(\Instr<13> ), .B(n141), .Y(\ExtImm<15> ) );
  NOR2BX1 U17 ( .AN(\Instr<14> ), .B(n141), .Y(\ExtImm<16> ) );
  NOR2X1 U18 ( .A(n141), .B(n143), .Y(\ExtImm<12> ) );
  NOR2X1 U19 ( .A(n141), .B(n142), .Y(\ExtImm<13> ) );
  NOR2BX1 U20 ( .AN(\Instr<12> ), .B(n141), .Y(\ExtImm<14> ) );
  NOR2BX1 U21 ( .AN(\Instr<15> ), .B(n155), .Y(\ExtImm<17> ) );
  NOR2BX1 U22 ( .AN(\Instr<16> ), .B(n155), .Y(\ExtImm<18> ) );
  NOR2BX1 U23 ( .AN(\Instr<18> ), .B(n155), .Y(\ExtImm<20> ) );
  NOR2BX1 U24 ( .AN(\Instr<20> ), .B(n155), .Y(\ExtImm<22> ) );
  NOR2BX1 U25 ( .AN(\Instr<17> ), .B(n155), .Y(\ExtImm<19> ) );
  NOR2BX1 U26 ( .AN(\Instr<19> ), .B(n155), .Y(\ExtImm<21> ) );
  INVX1 U27 ( .A(\Instr<2> ), .Y(n151) );
  INVX1 U28 ( .A(\Instr<3> ), .Y(n150) );
  INVX1 U29 ( .A(\Instr<0> ), .Y(n153) );
  INVX1 U30 ( .A(\Instr<1> ), .Y(n152) );
  NOR2BX1 U31 ( .AN(\Instr<22> ), .B(n141), .Y(\ExtImm<24> ) );
  NOR2BX1 U32 ( .AN(\Instr<21> ), .B(n141), .Y(\ExtImm<23> ) );
  INVX1 U33 ( .A(\ImmSrc<0> ), .Y(n154) );
  INVX1 U34 ( .A(\Instr<9> ), .Y(n144) );
  INVX1 U35 ( .A(\Instr<4> ), .Y(n149) );
  INVX1 U36 ( .A(\Instr<5> ), .Y(n148) );
  INVX1 U37 ( .A(\Instr<6> ), .Y(n147) );
  INVX1 U38 ( .A(\Instr<8> ), .Y(n145) );
  INVX1 U39 ( .A(\Instr<7> ), .Y(n146) );
  INVX1 U40 ( .A(\Instr<10> ), .Y(n143) );
  INVX1 U41 ( .A(\Instr<11> ), .Y(n142) );
  BUFX3 U42 ( .A(\ExtImm<25> ), .Y(\ExtImm<31> ) );
  BUFX3 U43 ( .A(\ExtImm<25> ), .Y(\ExtImm<30> ) );
  BUFX3 U44 ( .A(\ExtImm<25> ), .Y(\ExtImm<29> ) );
  BUFX3 U45 ( .A(\ExtImm<25> ), .Y(\ExtImm<28> ) );
  BUFX3 U46 ( .A(\ExtImm<25> ), .Y(\ExtImm<27> ) );
  BUFX3 U47 ( .A(\ExtImm<25> ), .Y(\ExtImm<26> ) );
  AND2X2 U48 ( .A(\Instr<23> ), .B(\ImmSrc<1> ), .Y(\ExtImm<25> ) );
endmodule


module alu_DW01_sub_0 ( .A({\A<31> , \A<30> , \A<29> , \A<28> , \A<27> , 
        \A<26> , \A<25> , \A<24> , \A<23> , \A<22> , \A<21> , \A<20> , \A<19> , 
        \A<18> , \A<17> , \A<16> , \A<15> , \A<14> , \A<13> , \A<12> , \A<11> , 
        \A<10> , \A<9> , \A<8> , \A<7> , \A<6> , \A<5> , \A<4> , \A<3> , 
        \A<2> , \A<1> , \A<0> }), .B({\B<31> , \B<30> , \B<29> , \B<28> , 
        \B<27> , \B<26> , \B<25> , \B<24> , \B<23> , \B<22> , \B<21> , \B<20> , 
        \B<19> , \B<18> , \B<17> , \B<16> , \B<15> , \B<14> , \B<13> , \B<12> , 
        \B<11> , \B<10> , \B<9> , \B<8> , \B<7> , \B<6> , \B<5> , \B<4> , 
        \B<3> , \B<2> , \B<1> , \B<0> }), CI, .DIFF({\DIFF<31> , \DIFF<30> , 
        \DIFF<29> , \DIFF<28> , \DIFF<27> , \DIFF<26> , \DIFF<25> , \DIFF<24> , 
        \DIFF<23> , \DIFF<22> , \DIFF<21> , \DIFF<20> , \DIFF<19> , \DIFF<18> , 
        \DIFF<17> , \DIFF<16> , \DIFF<15> , \DIFF<14> , \DIFF<13> , \DIFF<12> , 
        \DIFF<11> , \DIFF<10> , \DIFF<9> , \DIFF<8> , \DIFF<7> , \DIFF<6> , 
        \DIFF<5> , \DIFF<4> , \DIFF<3> , \DIFF<2> , \DIFF<1> , \DIFF<0> }), CO
 );
  input \A<31> , \A<30> , \A<29> , \A<28> , \A<27> , \A<26> , \A<25> , \A<24> ,
         \A<23> , \A<22> , \A<21> , \A<20> , \A<19> , \A<18> , \A<17> ,
         \A<16> , \A<15> , \A<14> , \A<13> , \A<12> , \A<11> , \A<10> , \A<9> ,
         \A<8> , \A<7> , \A<6> , \A<5> , \A<4> , \A<3> , \A<2> , \A<1> ,
         \A<0> , \B<31> , \B<30> , \B<29> , \B<28> , \B<27> , \B<26> , \B<25> ,
         \B<24> , \B<23> , \B<22> , \B<21> , \B<20> , \B<19> , \B<18> ,
         \B<17> , \B<16> , \B<15> , \B<14> , \B<13> , \B<12> , \B<11> ,
         \B<10> , \B<9> , \B<8> , \B<7> , \B<6> , \B<5> , \B<4> , \B<3> ,
         \B<2> , \B<1> , \B<0> , CI;
  output \DIFF<31> , \DIFF<30> , \DIFF<29> , \DIFF<28> , \DIFF<27> ,
         \DIFF<26> , \DIFF<25> , \DIFF<24> , \DIFF<23> , \DIFF<22> ,
         \DIFF<21> , \DIFF<20> , \DIFF<19> , \DIFF<18> , \DIFF<17> ,
         \DIFF<16> , \DIFF<15> , \DIFF<14> , \DIFF<13> , \DIFF<12> ,
         \DIFF<11> , \DIFF<10> , \DIFF<9> , \DIFF<8> , \DIFF<7> , \DIFF<6> ,
         \DIFF<5> , \DIFF<4> , \DIFF<3> , \DIFF<2> , \DIFF<1> , \DIFF<0> , CO;
  wire   \carry<31> , \carry<30> , \carry<29> , \carry<28> , \carry<27> ,
         \carry<26> , \carry<25> , \carry<24> , \carry<23> , \carry<22> ,
         \carry<21> , \carry<20> , \carry<19> , \carry<18> , \carry<17> ,
         \carry<16> , \carry<15> , \carry<14> , \carry<13> , \carry<12> ,
         \carry<11> , \carry<10> , \carry<9> , \carry<8> , \carry<7> ,
         \carry<6> , \carry<5> , \carry<4> , \carry<3> , \carry<2> ,
         \carry<1> , n187, n188, n189, n190, n191, n192, n193, n194, n195,
         n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206,
         n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217;

  ADDFX2 U2_29 ( .A(\A<29> ), .B(n188), .CI(\carry<29> ), .CO(\carry<30> ), 
        .S(\DIFF<29> ) );
  ADDFX2 U2_28 ( .A(\A<28> ), .B(n189), .CI(\carry<28> ), .CO(\carry<29> ), 
        .S(\DIFF<28> ) );
  ADDFX2 U2_27 ( .A(\A<27> ), .B(n190), .CI(\carry<27> ), .CO(\carry<28> ), 
        .S(\DIFF<27> ) );
  ADDFX2 U2_26 ( .A(\A<26> ), .B(n191), .CI(\carry<26> ), .CO(\carry<27> ), 
        .S(\DIFF<26> ) );
  ADDFX2 U2_25 ( .A(\A<25> ), .B(n192), .CI(\carry<25> ), .CO(\carry<26> ), 
        .S(\DIFF<25> ) );
  ADDFX2 U2_24 ( .A(\A<24> ), .B(n193), .CI(\carry<24> ), .CO(\carry<25> ), 
        .S(\DIFF<24> ) );
  ADDFX2 U2_23 ( .A(\A<23> ), .B(n194), .CI(\carry<23> ), .CO(\carry<24> ), 
        .S(\DIFF<23> ) );
  ADDFX2 U2_22 ( .A(\A<22> ), .B(n195), .CI(\carry<22> ), .CO(\carry<23> ), 
        .S(\DIFF<22> ) );
  ADDFX2 U2_21 ( .A(\A<21> ), .B(n196), .CI(\carry<21> ), .CO(\carry<22> ), 
        .S(\DIFF<21> ) );
  ADDFX2 U2_20 ( .A(\A<20> ), .B(n197), .CI(\carry<20> ), .CO(\carry<21> ), 
        .S(\DIFF<20> ) );
  ADDFX2 U2_19 ( .A(\A<19> ), .B(n198), .CI(\carry<19> ), .CO(\carry<20> ), 
        .S(\DIFF<19> ) );
  ADDFX2 U2_18 ( .A(\A<18> ), .B(n199), .CI(\carry<18> ), .CO(\carry<19> ), 
        .S(\DIFF<18> ) );
  ADDFX2 U2_17 ( .A(\A<17> ), .B(n200), .CI(\carry<17> ), .CO(\carry<18> ), 
        .S(\DIFF<17> ) );
  ADDFX2 U2_16 ( .A(\A<16> ), .B(n201), .CI(\carry<16> ), .CO(\carry<17> ), 
        .S(\DIFF<16> ) );
  ADDFX2 U2_15 ( .A(\A<15> ), .B(n202), .CI(\carry<15> ), .CO(\carry<16> ), 
        .S(\DIFF<15> ) );
  ADDFX2 U2_14 ( .A(\A<14> ), .B(n203), .CI(\carry<14> ), .CO(\carry<15> ), 
        .S(\DIFF<14> ) );
  ADDFX2 U2_13 ( .A(\A<13> ), .B(n204), .CI(\carry<13> ), .CO(\carry<14> ), 
        .S(\DIFF<13> ) );
  ADDFX2 U2_12 ( .A(\A<12> ), .B(n205), .CI(\carry<12> ), .CO(\carry<13> ), 
        .S(\DIFF<12> ) );
  ADDFX2 U2_11 ( .A(\A<11> ), .B(n206), .CI(\carry<11> ), .CO(\carry<12> ), 
        .S(\DIFF<11> ) );
  ADDFX2 U2_10 ( .A(\A<10> ), .B(n207), .CI(\carry<10> ), .CO(\carry<11> ), 
        .S(\DIFF<10> ) );
  ADDFX2 U2_9 ( .A(\A<9> ), .B(n208), .CI(\carry<9> ), .CO(\carry<10> ), .S(
        \DIFF<9> ) );
  ADDFX2 U2_8 ( .A(\A<8> ), .B(n209), .CI(\carry<8> ), .CO(\carry<9> ), .S(
        \DIFF<8> ) );
  ADDFX2 U2_7 ( .A(\A<7> ), .B(n210), .CI(\carry<7> ), .CO(\carry<8> ), .S(
        \DIFF<7> ) );
  ADDFX2 U2_6 ( .A(\A<6> ), .B(n211), .CI(\carry<6> ), .CO(\carry<7> ), .S(
        \DIFF<6> ) );
  ADDFX2 U2_5 ( .A(\A<5> ), .B(n212), .CI(\carry<5> ), .CO(\carry<6> ), .S(
        \DIFF<5> ) );
  ADDFX2 U2_4 ( .A(\A<4> ), .B(n213), .CI(\carry<4> ), .CO(\carry<5> ), .S(
        \DIFF<4> ) );
  ADDFX2 U2_3 ( .A(\A<3> ), .B(n214), .CI(\carry<3> ), .CO(\carry<4> ), .S(
        \DIFF<3> ) );
  ADDFX2 U2_2 ( .A(\A<2> ), .B(n215), .CI(\carry<2> ), .CO(\carry<3> ), .S(
        \DIFF<2> ) );
  ADDFX2 U2_1 ( .A(\A<1> ), .B(n216), .CI(\carry<1> ), .CO(\carry<2> ), .S(
        \DIFF<1> ) );
  ADDFX2 U2_30 ( .A(\A<30> ), .B(n187), .CI(\carry<30> ), .CO(\carry<31> ), 
        .S(\DIFF<30> ) );
  XNOR3X2 U1 ( .A(\A<31> ), .B(\B<31> ), .C(\carry<31> ), .Y(\DIFF<31> ) );
  INVX1 U2 ( .A(\B<0> ), .Y(n217) );
  INVX1 U3 ( .A(\B<30> ), .Y(n187) );
  INVX1 U4 ( .A(\B<1> ), .Y(n216) );
  OR2X2 U5 ( .A(\A<0> ), .B(n217), .Y(\carry<1> ) );
  INVX1 U6 ( .A(\B<2> ), .Y(n215) );
  INVX1 U7 ( .A(\B<3> ), .Y(n214) );
  INVX1 U8 ( .A(\B<4> ), .Y(n213) );
  INVX1 U9 ( .A(\B<5> ), .Y(n212) );
  INVX1 U10 ( .A(\B<6> ), .Y(n211) );
  INVX1 U11 ( .A(\B<7> ), .Y(n210) );
  INVX1 U12 ( .A(\B<8> ), .Y(n209) );
  INVX1 U13 ( .A(\B<9> ), .Y(n208) );
  INVX1 U14 ( .A(\B<10> ), .Y(n207) );
  INVX1 U15 ( .A(\B<11> ), .Y(n206) );
  INVX1 U16 ( .A(\B<12> ), .Y(n205) );
  INVX1 U17 ( .A(\B<13> ), .Y(n204) );
  INVX1 U18 ( .A(\B<14> ), .Y(n203) );
  INVX1 U19 ( .A(\B<15> ), .Y(n202) );
  INVX1 U20 ( .A(\B<16> ), .Y(n201) );
  INVX1 U21 ( .A(\B<17> ), .Y(n200) );
  INVX1 U22 ( .A(\B<18> ), .Y(n199) );
  INVX1 U23 ( .A(\B<19> ), .Y(n198) );
  INVX1 U24 ( .A(\B<20> ), .Y(n197) );
  INVX1 U25 ( .A(\B<21> ), .Y(n196) );
  INVX1 U26 ( .A(\B<22> ), .Y(n195) );
  INVX1 U27 ( .A(\B<23> ), .Y(n194) );
  INVX1 U28 ( .A(\B<24> ), .Y(n193) );
  INVX1 U29 ( .A(\B<25> ), .Y(n192) );
  INVX1 U30 ( .A(\B<26> ), .Y(n191) );
  INVX1 U31 ( .A(\B<27> ), .Y(n190) );
  INVX1 U32 ( .A(\B<28> ), .Y(n189) );
  INVX1 U33 ( .A(\B<29> ), .Y(n188) );
  XNOR2X1 U34 ( .A(n217), .B(\A<0> ), .Y(\DIFF<0> ) );
endmodule


module alu_DW01_add_0 ( .A({\A<32> , \A<31> , \A<30> , \A<29> , \A<28> , 
        \A<27> , \A<26> , \A<25> , \A<24> , \A<23> , \A<22> , \A<21> , \A<20> , 
        \A<19> , \A<18> , \A<17> , \A<16> , \A<15> , \A<14> , \A<13> , \A<12> , 
        \A<11> , \A<10> , \A<9> , \A<8> , \A<7> , \A<6> , \A<5> , \A<4> , 
        \A<3> , \A<2> , \A<1> , \A<0> }), .B({\B<32> , \B<31> , \B<30> , 
        \B<29> , \B<28> , \B<27> , \B<26> , \B<25> , \B<24> , \B<23> , \B<22> , 
        \B<21> , \B<20> , \B<19> , \B<18> , \B<17> , \B<16> , \B<15> , \B<14> , 
        \B<13> , \B<12> , \B<11> , \B<10> , \B<9> , \B<8> , \B<7> , \B<6> , 
        \B<5> , \B<4> , \B<3> , \B<2> , \B<1> , \B<0> }), CI, .SUM({\SUM<32> , 
        \SUM<31> , \SUM<30> , \SUM<29> , \SUM<28> , \SUM<27> , \SUM<26> , 
        \SUM<25> , \SUM<24> , \SUM<23> , \SUM<22> , \SUM<21> , \SUM<20> , 
        \SUM<19> , \SUM<18> , \SUM<17> , \SUM<16> , \SUM<15> , \SUM<14> , 
        \SUM<13> , \SUM<12> , \SUM<11> , \SUM<10> , \SUM<9> , \SUM<8> , 
        \SUM<7> , \SUM<6> , \SUM<5> , \SUM<4> , \SUM<3> , \SUM<2> , \SUM<1> , 
        \SUM<0> }), CO );
  input \A<32> , \A<31> , \A<30> , \A<29> , \A<28> , \A<27> , \A<26> , \A<25> ,
         \A<24> , \A<23> , \A<22> , \A<21> , \A<20> , \A<19> , \A<18> ,
         \A<17> , \A<16> , \A<15> , \A<14> , \A<13> , \A<12> , \A<11> ,
         \A<10> , \A<9> , \A<8> , \A<7> , \A<6> , \A<5> , \A<4> , \A<3> ,
         \A<2> , \A<1> , \A<0> , \B<32> , \B<31> , \B<30> , \B<29> , \B<28> ,
         \B<27> , \B<26> , \B<25> , \B<24> , \B<23> , \B<22> , \B<21> ,
         \B<20> , \B<19> , \B<18> , \B<17> , \B<16> , \B<15> , \B<14> ,
         \B<13> , \B<12> , \B<11> , \B<10> , \B<9> , \B<8> , \B<7> , \B<6> ,
         \B<5> , \B<4> , \B<3> , \B<2> , \B<1> , \B<0> , CI;
  output \SUM<32> , \SUM<31> , \SUM<30> , \SUM<29> , \SUM<28> , \SUM<27> ,
         \SUM<26> , \SUM<25> , \SUM<24> , \SUM<23> , \SUM<22> , \SUM<21> ,
         \SUM<20> , \SUM<19> , \SUM<18> , \SUM<17> , \SUM<16> , \SUM<15> ,
         \SUM<14> , \SUM<13> , \SUM<12> , \SUM<11> , \SUM<10> , \SUM<9> ,
         \SUM<8> , \SUM<7> , \SUM<6> , \SUM<5> , \SUM<4> , \SUM<3> , \SUM<2> ,
         \SUM<1> , \SUM<0> , CO;
  wire   \carry<31> , \carry<30> , \carry<29> , \carry<28> , \carry<27> ,
         \carry<26> , \carry<25> , \carry<24> , \carry<23> , \carry<22> ,
         \carry<21> , \carry<20> , \carry<19> , \carry<18> , \carry<17> ,
         \carry<16> , \carry<15> , \carry<14> , \carry<13> , \carry<12> ,
         \carry<11> , \carry<10> , \carry<9> , \carry<8> , \carry<7> ,
         \carry<6> , \carry<5> , \carry<4> , \carry<3> , \carry<2> ,
         \carry<1> ;

  ADDFX2 U1_30 ( .A(\A<30> ), .B(\B<30> ), .CI(\carry<30> ), .CO(\carry<31> ), 
        .S(\SUM<30> ) );
  ADDFX2 U1_29 ( .A(\A<29> ), .B(\B<29> ), .CI(\carry<29> ), .CO(\carry<30> ), 
        .S(\SUM<29> ) );
  ADDFX2 U1_28 ( .A(\A<28> ), .B(\B<28> ), .CI(\carry<28> ), .CO(\carry<29> ), 
        .S(\SUM<28> ) );
  ADDFX2 U1_27 ( .A(\A<27> ), .B(\B<27> ), .CI(\carry<27> ), .CO(\carry<28> ), 
        .S(\SUM<27> ) );
  ADDFX2 U1_26 ( .A(\A<26> ), .B(\B<26> ), .CI(\carry<26> ), .CO(\carry<27> ), 
        .S(\SUM<26> ) );
  ADDFX2 U1_25 ( .A(\A<25> ), .B(\B<25> ), .CI(\carry<25> ), .CO(\carry<26> ), 
        .S(\SUM<25> ) );
  ADDFX2 U1_24 ( .A(\A<24> ), .B(\B<24> ), .CI(\carry<24> ), .CO(\carry<25> ), 
        .S(\SUM<24> ) );
  ADDFX2 U1_23 ( .A(\A<23> ), .B(\B<23> ), .CI(\carry<23> ), .CO(\carry<24> ), 
        .S(\SUM<23> ) );
  ADDFX2 U1_22 ( .A(\A<22> ), .B(\B<22> ), .CI(\carry<22> ), .CO(\carry<23> ), 
        .S(\SUM<22> ) );
  ADDFX2 U1_21 ( .A(\A<21> ), .B(\B<21> ), .CI(\carry<21> ), .CO(\carry<22> ), 
        .S(\SUM<21> ) );
  ADDFX2 U1_20 ( .A(\A<20> ), .B(\B<20> ), .CI(\carry<20> ), .CO(\carry<21> ), 
        .S(\SUM<20> ) );
  ADDFX2 U1_19 ( .A(\A<19> ), .B(\B<19> ), .CI(\carry<19> ), .CO(\carry<20> ), 
        .S(\SUM<19> ) );
  ADDFX2 U1_18 ( .A(\A<18> ), .B(\B<18> ), .CI(\carry<18> ), .CO(\carry<19> ), 
        .S(\SUM<18> ) );
  ADDFX2 U1_17 ( .A(\A<17> ), .B(\B<17> ), .CI(\carry<17> ), .CO(\carry<18> ), 
        .S(\SUM<17> ) );
  ADDFX2 U1_16 ( .A(\A<16> ), .B(\B<16> ), .CI(\carry<16> ), .CO(\carry<17> ), 
        .S(\SUM<16> ) );
  ADDFX2 U1_15 ( .A(\A<15> ), .B(\B<15> ), .CI(\carry<15> ), .CO(\carry<16> ), 
        .S(\SUM<15> ) );
  ADDFX2 U1_14 ( .A(\A<14> ), .B(\B<14> ), .CI(\carry<14> ), .CO(\carry<15> ), 
        .S(\SUM<14> ) );
  ADDFX2 U1_13 ( .A(\A<13> ), .B(\B<13> ), .CI(\carry<13> ), .CO(\carry<14> ), 
        .S(\SUM<13> ) );
  ADDFX2 U1_12 ( .A(\A<12> ), .B(\B<12> ), .CI(\carry<12> ), .CO(\carry<13> ), 
        .S(\SUM<12> ) );
  ADDFX2 U1_9 ( .A(\A<9> ), .B(\B<9> ), .CI(\carry<9> ), .CO(\carry<10> ), .S(
        \SUM<9> ) );
  ADDFX2 U1_11 ( .A(\A<11> ), .B(\B<11> ), .CI(\carry<11> ), .CO(\carry<12> ), 
        .S(\SUM<11> ) );
  ADDFX2 U1_10 ( .A(\A<10> ), .B(\B<10> ), .CI(\carry<10> ), .CO(\carry<11> ), 
        .S(\SUM<10> ) );
  ADDFX2 U1_8 ( .A(\A<8> ), .B(\B<8> ), .CI(\carry<8> ), .CO(\carry<9> ), .S(
        \SUM<8> ) );
  ADDFX2 U1_7 ( .A(\A<7> ), .B(\B<7> ), .CI(\carry<7> ), .CO(\carry<8> ), .S(
        \SUM<7> ) );
  ADDFX2 U1_6 ( .A(\A<6> ), .B(\B<6> ), .CI(\carry<6> ), .CO(\carry<7> ), .S(
        \SUM<6> ) );
  ADDFX2 U1_5 ( .A(\A<5> ), .B(\B<5> ), .CI(\carry<5> ), .CO(\carry<6> ), .S(
        \SUM<5> ) );
  ADDFX2 U1_4 ( .A(\A<4> ), .B(\B<4> ), .CI(\carry<4> ), .CO(\carry<5> ), .S(
        \SUM<4> ) );
  ADDFX2 U1_3 ( .A(\A<3> ), .B(\B<3> ), .CI(\carry<3> ), .CO(\carry<4> ), .S(
        \SUM<3> ) );
  ADDFX2 U1_2 ( .A(\A<2> ), .B(\B<2> ), .CI(\carry<2> ), .CO(\carry<3> ), .S(
        \SUM<2> ) );
  ADDFX2 U1_1 ( .A(\A<1> ), .B(\B<1> ), .CI(\carry<1> ), .CO(\carry<2> ), .S(
        \SUM<1> ) );
  ADDFX2 U1_31 ( .A(\A<31> ), .B(\B<31> ), .CI(\carry<31> ), .CO(\SUM<32> ), 
        .S(\SUM<31> ) );
  AND2X2 U1 ( .A(\B<0> ), .B(\A<0> ), .Y(\carry<1> ) );
  XOR2X1 U2 ( .A(\B<0> ), .B(\A<0> ), .Y(\SUM<0> ) );
endmodule


module alu ( .a({\a<31> , \a<30> , \a<29> , \a<28> , \a<27> , \a<26> , \a<25> , 
        \a<24> , \a<23> , \a<22> , \a<21> , \a<20> , \a<19> , \a<18> , \a<17> , 
        \a<16> , \a<15> , \a<14> , \a<13> , \a<12> , \a<11> , \a<10> , \a<9> , 
        \a<8> , \a<7> , \a<6> , \a<5> , \a<4> , \a<3> , \a<2> , \a<1> , \a<0> 
        }), .b({\b<31> , \b<30> , \b<29> , \b<28> , \b<27> , \b<26> , \b<25> , 
        \b<24> , \b<23> , \b<22> , \b<21> , \b<20> , \b<19> , \b<18> , \b<17> , 
        \b<16> , \b<15> , \b<14> , \b<13> , \b<12> , \b<11> , \b<10> , \b<9> , 
        \b<8> , \b<7> , \b<6> , \b<5> , \b<4> , \b<3> , \b<2> , \b<1> , \b<0> 
        }), .ALUControl({\ALUControl<1> , \ALUControl<0> }), .Result({
        \Result<31> , \Result<30> , \Result<29> , \Result<28> , \Result<27> , 
        \Result<26> , \Result<25> , \Result<24> , \Result<23> , \Result<22> , 
        \Result<21> , \Result<20> , \Result<19> , \Result<18> , \Result<17> , 
        \Result<16> , \Result<15> , \Result<14> , \Result<13> , \Result<12> , 
        \Result<11> , \Result<10> , \Result<9> , \Result<8> , \Result<7> , 
        \Result<6> , \Result<5> , \Result<4> , \Result<3> , \Result<2> , 
        \Result<1> , \Result<0> }), .ALUFlags({\ALUFlags<3> , \ALUFlags<2> , 
        \ALUFlags<1> , \ALUFlags<0> }) );
  input \a<31> , \a<30> , \a<29> , \a<28> , \a<27> , \a<26> , \a<25> , \a<24> ,
         \a<23> , \a<22> , \a<21> , \a<20> , \a<19> , \a<18> , \a<17> ,
         \a<16> , \a<15> , \a<14> , \a<13> , \a<12> , \a<11> , \a<10> , \a<9> ,
         \a<8> , \a<7> , \a<6> , \a<5> , \a<4> , \a<3> , \a<2> , \a<1> ,
         \a<0> , \b<31> , \b<30> , \b<29> , \b<28> , \b<27> , \b<26> , \b<25> ,
         \b<24> , \b<23> , \b<22> , \b<21> , \b<20> , \b<19> , \b<18> ,
         \b<17> , \b<16> , \b<15> , \b<14> , \b<13> , \b<12> , \b<11> ,
         \b<10> , \b<9> , \b<8> , \b<7> , \b<6> , \b<5> , \b<4> , \b<3> ,
         \b<2> , \b<1> , \b<0> , \ALUControl<1> , \ALUControl<0> ;
  output \Result<31> , \Result<30> , \Result<29> , \Result<28> , \Result<27> ,
         \Result<26> , \Result<25> , \Result<24> , \Result<23> , \Result<22> ,
         \Result<21> , \Result<20> , \Result<19> , \Result<18> , \Result<17> ,
         \Result<16> , \Result<15> , \Result<14> , \Result<13> , \Result<12> ,
         \Result<11> , \Result<10> , \Result<9> , \Result<8> , \Result<7> ,
         \Result<6> , \Result<5> , \Result<4> , \Result<3> , \Result<2> ,
         \Result<1> , \Result<0> , \ALUFlags<3> , \ALUFlags<2> , \ALUFlags<1> ,
         \ALUFlags<0> ;
  wire   N13, N14, N15, N16, N17, N18, N19, N20, N21, N22, N23, N24, N25, N26,
         N27, N28, N29, N30, N31, N32, N33, N34, N35, N36, N37, N38, N39, N40,
         N41, N42, N43, N44, N45, N46, N47, N48, N49, N50, N51, N52, N53, N54,
         N55, N56, N57, N58, N59, N60, N61, N62, N63, N64, N65, N66, N67, N68,
         N69, N70, N71, N72, N73, N74, N75, N76, N77, N173, n6, n7, n8, n9,
         n10, n11, n12, n13, n14, n17, n18, n19, n20, n21, n22, n23, n24, n25,
         n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39,
         n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53,
         n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67,
         n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81,
         n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95,
         n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107,
         n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n225,
         n226, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237,
         n238, n239, n240, n241, n242;
  assign \ALUFlags<2>  = N173;

  alu_DW01_sub_0 sub_466 ( .A({\a<31> , \a<30> , \a<29> , \a<28> , \a<27> , 
        \a<26> , \a<25> , \a<24> , \a<23> , \a<22> , \a<21> , \a<20> , \a<19> , 
        \a<18> , \a<17> , \a<16> , \a<15> , \a<14> , \a<13> , \a<12> , \a<11> , 
        \a<10> , \a<9> , \a<8> , \a<7> , \a<6> , \a<5> , \a<4> , \a<3> , 
        \a<2> , \a<1> , \a<0> }), .B({\b<31> , \b<30> , \b<29> , \b<28> , 
        \b<27> , \b<26> , \b<25> , \b<24> , \b<23> , \b<22> , \b<21> , \b<20> , 
        \b<19> , \b<18> , \b<17> , \b<16> , \b<15> , \b<14> , \b<13> , \b<12> , 
        \b<11> , \b<10> , \b<9> , \b<8> , \b<7> , \b<6> , \b<5> , \b<4> , 
        \b<3> , \b<2> , \b<1> , \b<0> }), .CI(1'b0), .DIFF({N77, N76, N75, N74, 
        N73, N72, N71, N70, N69, N68, N67, N66, N65, N64, N63, N62, N61, N60, 
        N59, N58, N57, N56, N55, N54, N53, N52, N51, N50, N49, N48, N47, N46})
         );
  alu_DW01_add_0 add_465 ( .A({1'b0, \a<31> , \a<30> , \a<29> , \a<28> , 
        \a<27> , \a<26> , \a<25> , \a<24> , \a<23> , \a<22> , \a<21> , \a<20> , 
        \a<19> , \a<18> , \a<17> , \a<16> , \a<15> , \a<14> , \a<13> , \a<12> , 
        \a<11> , \a<10> , \a<9> , \a<8> , \a<7> , \a<6> , \a<5> , \a<4> , 
        \a<3> , \a<2> , \a<1> , \a<0> }), .B({1'b0, \b<31> , \b<30> , \b<29> , 
        \b<28> , \b<27> , \b<26> , \b<25> , \b<24> , \b<23> , \b<22> , \b<21> , 
        \b<20> , \b<19> , \b<18> , \b<17> , \b<16> , \b<15> , \b<14> , \b<13> , 
        \b<12> , \b<11> , \b<10> , \b<9> , \b<8> , \b<7> , \b<6> , \b<5> , 
        \b<4> , \b<3> , \b<2> , \b<1> , \b<0> }), .CI(1'b0), .SUM({N45, N44, 
        N43, N42, N41, N40, N39, N38, N37, N36, N35, N34, N33, N32, N31, N30, 
        N29, N28, N27, N26, N25, N24, N23, N22, N21, N20, N19, N18, N17, N16, 
        N15, N14, N13}) );
  OR2X2 U4 ( .A(n240), .B(\ALUControl<0> ), .Y(n225) );
  CLKINVX3 U5 ( .A(n231), .Y(n232) );
  INVX1 U6 ( .A(n226), .Y(n234) );
  INVX1 U7 ( .A(n226), .Y(n233) );
  INVX1 U8 ( .A(n237), .Y(n236) );
  INVX1 U9 ( .A(n226), .Y(n235) );
  CLKINVX3 U10 ( .A(n242), .Y(n241) );
  CLKINVX3 U11 ( .A(n242), .Y(n240) );
  INVX1 U12 ( .A(\ALUControl<1> ), .Y(n242) );
  CLKINVX3 U13 ( .A(n230), .Y(n229) );
  CLKINVX3 U14 ( .A(n225), .Y(n238) );
  CLKINVX3 U15 ( .A(n225), .Y(n239) );
  INVX1 U16 ( .A(n231), .Y(n237) );
  OR4X2 U17 ( .A(\Result<31> ), .B(\Result<3> ), .C(\Result<4> ), .D(
        \Result<5> ), .Y(n66) );
  OR4X2 U18 ( .A(n63), .B(n64), .C(n65), .D(n66), .Y(n6) );
  OR4X2 U19 ( .A(\Result<6> ), .B(\Result<7> ), .C(\Result<8> ), .D(
        \Result<9> ), .Y(n65) );
  OR4X2 U20 ( .A(\Result<24> ), .B(\Result<25> ), .C(\Result<26> ), .D(
        \Result<27> ), .Y(n64) );
  OR4X2 U21 ( .A(\Result<28> ), .B(\Result<29> ), .C(\Result<2> ), .D(
        \Result<30> ), .Y(n63) );
  OR4X2 U22 ( .A(\Result<20> ), .B(\Result<21> ), .C(\Result<22> ), .D(
        \Result<23> ), .Y(n10) );
  OR4X2 U23 ( .A(\Result<17> ), .B(\Result<18> ), .C(\Result<19> ), .D(
        \Result<1> ), .Y(n11) );
  OR4X2 U24 ( .A(\Result<0> ), .B(\Result<10> ), .C(\Result<11> ), .D(
        \Result<12> ), .Y(n9) );
  OR4X2 U25 ( .A(\Result<13> ), .B(\Result<14> ), .C(\Result<15> ), .D(
        \Result<16> ), .Y(n8) );
  INVX1 U26 ( .A(n226), .Y(n231) );
  CLKINVX3 U27 ( .A(n230), .Y(n228) );
  INVX1 U28 ( .A(n17), .Y(n230) );
  AOI22X1 U29 ( .A0(N77), .A1(n228), .B0(\a<31> ), .B1(n237), .Y(n115) );
  AOI22X1 U30 ( .A0(\b<31> ), .A1(n117), .B0(N44), .B1(n239), .Y(n116) );
  NAND2X1 U31 ( .A(n88), .B(n89), .Y(\Result<27> ) );
  AOI22X1 U32 ( .A0(N73), .A1(n228), .B0(\a<27> ), .B1(n232), .Y(n88) );
  AOI22X1 U33 ( .A0(\b<27> ), .A1(n90), .B0(N40), .B1(n239), .Y(n89) );
  OAI2BB1X1 U34 ( .A0N(n241), .A1N(\a<27> ), .B0(n235), .Y(n90) );
  NAND2X1 U35 ( .A(n106), .B(n107), .Y(\Result<29> ) );
  AOI22X1 U36 ( .A0(N75), .A1(n228), .B0(\a<29> ), .B1(n226), .Y(n106) );
  AOI22X1 U37 ( .A0(\b<29> ), .A1(n108), .B0(N42), .B1(n239), .Y(n107) );
  OAI2BB1X1 U38 ( .A0N(n241), .A1N(\a<29> ), .B0(n231), .Y(n108) );
  NAND2X1 U39 ( .A(n91), .B(n92), .Y(\Result<26> ) );
  AOI22X1 U40 ( .A0(N72), .A1(n228), .B0(\a<26> ), .B1(n232), .Y(n91) );
  AOI22X1 U41 ( .A0(\b<26> ), .A1(n93), .B0(N39), .B1(n239), .Y(n92) );
  OAI2BB1X1 U42 ( .A0N(n241), .A1N(\a<26> ), .B0(n236), .Y(n93) );
  NAND2X1 U43 ( .A(n109), .B(n110), .Y(\Result<28> ) );
  AOI22X1 U44 ( .A0(N74), .A1(n228), .B0(\a<28> ), .B1(n226), .Y(n109) );
  AOI22X1 U45 ( .A0(\b<28> ), .A1(n111), .B0(N41), .B1(n239), .Y(n110) );
  OAI2BB1X1 U46 ( .A0N(n241), .A1N(\a<28> ), .B0(n236), .Y(n111) );
  NAND2X1 U47 ( .A(n100), .B(n101), .Y(\Result<30> ) );
  AOI22X1 U48 ( .A0(N76), .A1(n228), .B0(\a<30> ), .B1(n226), .Y(n100) );
  AOI22X1 U49 ( .A0(\b<30> ), .A1(n102), .B0(N43), .B1(n239), .Y(n101) );
  OAI2BB1X1 U50 ( .A0N(n241), .A1N(\a<30> ), .B0(n231), .Y(n102) );
  NAND2X1 U51 ( .A(n30), .B(n31), .Y(\Result<22> ) );
  AOI22X1 U52 ( .A0(N68), .A1(n228), .B0(\a<22> ), .B1(n232), .Y(n30) );
  AOI22X1 U53 ( .A0(\b<22> ), .A1(n32), .B0(N35), .B1(n239), .Y(n31) );
  OAI2BB1X1 U54 ( .A0N(n240), .A1N(\a<22> ), .B0(n234), .Y(n32) );
  NAND2X1 U55 ( .A(n33), .B(n34), .Y(\Result<21> ) );
  AOI22X1 U56 ( .A0(N67), .A1(n228), .B0(\a<21> ), .B1(n237), .Y(n33) );
  AOI22X1 U57 ( .A0(\b<21> ), .A1(n35), .B0(N34), .B1(n239), .Y(n34) );
  OAI2BB1X1 U58 ( .A0N(n240), .A1N(\a<21> ), .B0(n235), .Y(n35) );
  NAND2X1 U59 ( .A(n94), .B(n95), .Y(\Result<25> ) );
  AOI22X1 U60 ( .A0(N71), .A1(n228), .B0(\a<25> ), .B1(n232), .Y(n94) );
  AOI22X1 U61 ( .A0(\b<25> ), .A1(n96), .B0(N38), .B1(n239), .Y(n95) );
  OAI2BB1X1 U62 ( .A0N(n241), .A1N(\a<25> ), .B0(n236), .Y(n96) );
  NAND2X1 U63 ( .A(n27), .B(n28), .Y(\Result<23> ) );
  AOI22X1 U64 ( .A0(N69), .A1(n228), .B0(\a<23> ), .B1(n237), .Y(n27) );
  AOI22X1 U65 ( .A0(\b<23> ), .A1(n29), .B0(N36), .B1(n239), .Y(n28) );
  OAI2BB1X1 U66 ( .A0N(n240), .A1N(\a<23> ), .B0(n235), .Y(n29) );
  NAND2X1 U67 ( .A(n97), .B(n98), .Y(\Result<24> ) );
  AOI22X1 U68 ( .A0(N70), .A1(n228), .B0(\a<24> ), .B1(n226), .Y(n97) );
  AOI22X1 U69 ( .A0(\b<24> ), .A1(n99), .B0(N37), .B1(n239), .Y(n98) );
  OAI2BB1X1 U70 ( .A0N(n241), .A1N(\a<24> ), .B0(n231), .Y(n99) );
  XNOR2X1 U71 ( .A(\a<31> ), .B(\Result<31> ), .Y(n112) );
  NAND2X1 U72 ( .A(n18), .B(n19), .Y(\Result<19> ) );
  AOI22X1 U73 ( .A0(N65), .A1(n228), .B0(\a<19> ), .B1(n237), .Y(n18) );
  AOI22X1 U74 ( .A0(\b<19> ), .A1(n20), .B0(N32), .B1(n239), .Y(n19) );
  OAI2BB1X1 U75 ( .A0N(n240), .A1N(\a<19> ), .B0(n236), .Y(n20) );
  NAND2X1 U76 ( .A(n21), .B(n22), .Y(\Result<18> ) );
  AOI22X1 U77 ( .A0(N64), .A1(n228), .B0(\a<18> ), .B1(n237), .Y(n21) );
  AOI22X1 U78 ( .A0(\b<18> ), .A1(n23), .B0(N31), .B1(n239), .Y(n22) );
  OAI2BB1X1 U79 ( .A0N(n240), .A1N(\a<18> ), .B0(n235), .Y(n23) );
  NAND2X1 U80 ( .A(n24), .B(n25), .Y(\Result<17> ) );
  AOI22X1 U81 ( .A0(N63), .A1(n228), .B0(\a<17> ), .B1(n232), .Y(n24) );
  AOI22X1 U82 ( .A0(\b<17> ), .A1(n26), .B0(N30), .B1(n239), .Y(n25) );
  OAI2BB1X1 U83 ( .A0N(n240), .A1N(\a<17> ), .B0(n234), .Y(n26) );
  NAND2X1 U84 ( .A(n36), .B(n37), .Y(\Result<20> ) );
  AOI22X1 U85 ( .A0(N66), .A1(n228), .B0(\a<20> ), .B1(n232), .Y(n36) );
  AOI22X1 U86 ( .A0(\b<20> ), .A1(n38), .B0(N33), .B1(n239), .Y(n37) );
  OAI2BB1X1 U87 ( .A0N(n240), .A1N(\a<20> ), .B0(n234), .Y(n38) );
  NAND2X1 U88 ( .A(n39), .B(n40), .Y(\Result<12> ) );
  AOI22X1 U89 ( .A0(N58), .A1(n229), .B0(\a<12> ), .B1(n232), .Y(n39) );
  AOI22X1 U90 ( .A0(\b<12> ), .A1(n41), .B0(N25), .B1(n239), .Y(n40) );
  OAI2BB1X1 U91 ( .A0N(n240), .A1N(\a<12> ), .B0(n234), .Y(n41) );
  NAND2X1 U92 ( .A(n54), .B(n55), .Y(\Result<15> ) );
  AOI22X1 U93 ( .A0(N61), .A1(n229), .B0(\a<15> ), .B1(n232), .Y(n54) );
  AOI22X1 U94 ( .A0(\b<15> ), .A1(n56), .B0(N28), .B1(n238), .Y(n55) );
  OAI2BB1X1 U95 ( .A0N(n241), .A1N(\a<15> ), .B0(n231), .Y(n56) );
  NAND2X1 U96 ( .A(n57), .B(n58), .Y(\Result<14> ) );
  AOI22X1 U97 ( .A0(N60), .A1(n229), .B0(\a<14> ), .B1(n232), .Y(n57) );
  AOI22X1 U98 ( .A0(\b<14> ), .A1(n59), .B0(N27), .B1(n238), .Y(n58) );
  OAI2BB1X1 U99 ( .A0N(n241), .A1N(\a<14> ), .B0(n233), .Y(n59) );
  NAND2X1 U100 ( .A(n60), .B(n61), .Y(\Result<13> ) );
  AOI22X1 U101 ( .A0(N59), .A1(n229), .B0(\a<13> ), .B1(n232), .Y(n60) );
  AOI22X1 U102 ( .A0(\b<13> ), .A1(n62), .B0(N26), .B1(n238), .Y(n61) );
  OAI2BB1X1 U103 ( .A0N(n241), .A1N(\a<13> ), .B0(n234), .Y(n62) );
  NAND2X1 U104 ( .A(n51), .B(n52), .Y(\Result<16> ) );
  AOI22X1 U105 ( .A0(N62), .A1(n229), .B0(\a<16> ), .B1(n232), .Y(n51) );
  AOI22X1 U106 ( .A0(\b<16> ), .A1(n53), .B0(N29), .B1(n238), .Y(n52) );
  OAI2BB1X1 U107 ( .A0N(n241), .A1N(\a<16> ), .B0(n233), .Y(n53) );
  NAND2X1 U108 ( .A(n79), .B(n80), .Y(\Result<8> ) );
  AOI22X1 U109 ( .A0(N54), .A1(n228), .B0(\a<8> ), .B1(n232), .Y(n79) );
  AOI22X1 U110 ( .A0(\b<8> ), .A1(n81), .B0(N21), .B1(n238), .Y(n80) );
  OAI2BB1X1 U111 ( .A0N(n241), .A1N(\a<8> ), .B0(n234), .Y(n81) );
  NAND2X1 U112 ( .A(n42), .B(n43), .Y(\Result<11> ) );
  AOI22X1 U113 ( .A0(N57), .A1(n229), .B0(\a<11> ), .B1(n232), .Y(n42) );
  AOI22X1 U114 ( .A0(\b<11> ), .A1(n44), .B0(N24), .B1(n239), .Y(n43) );
  OAI2BB1X1 U115 ( .A0N(n240), .A1N(\a<11> ), .B0(n236), .Y(n44) );
  NAND2X1 U116 ( .A(n82), .B(n83), .Y(\Result<7> ) );
  AOI22X1 U117 ( .A0(N53), .A1(n228), .B0(\a<7> ), .B1(n232), .Y(n82) );
  AOI22X1 U118 ( .A0(\b<7> ), .A1(n84), .B0(N20), .B1(n238), .Y(n83) );
  OAI2BB1X1 U119 ( .A0N(n241), .A1N(\a<7> ), .B0(n234), .Y(n84) );
  NAND2X1 U120 ( .A(n45), .B(n46), .Y(\Result<10> ) );
  AOI22X1 U121 ( .A0(N56), .A1(n229), .B0(\a<10> ), .B1(n232), .Y(n45) );
  AOI22X1 U122 ( .A0(\b<10> ), .A1(n47), .B0(N23), .B1(n239), .Y(n46) );
  OAI2BB1X1 U123 ( .A0N(n241), .A1N(\a<10> ), .B0(n236), .Y(n47) );
  NAND2X1 U124 ( .A(n76), .B(n77), .Y(\Result<9> ) );
  AOI22X1 U125 ( .A0(N55), .A1(n229), .B0(n232), .B1(\a<9> ), .Y(n76) );
  AOI22X1 U126 ( .A0(\b<9> ), .A1(n78), .B0(N22), .B1(n238), .Y(n77) );
  OAI2BB1X1 U127 ( .A0N(n241), .A1N(\a<9> ), .B0(n233), .Y(n78) );
  NAND2X1 U128 ( .A(n103), .B(n104), .Y(\Result<2> ) );
  AOI22X1 U129 ( .A0(N48), .A1(n228), .B0(\a<2> ), .B1(n237), .Y(n103) );
  AOI22X1 U130 ( .A0(\b<2> ), .A1(n105), .B0(N15), .B1(n239), .Y(n104) );
  OAI2BB1X1 U131 ( .A0N(n241), .A1N(\a<2> ), .B0(n233), .Y(n105) );
  NAND2X1 U132 ( .A(n70), .B(n71), .Y(\Result<4> ) );
  AOI22X1 U133 ( .A0(N50), .A1(n229), .B0(\a<4> ), .B1(n232), .Y(n70) );
  AOI22X1 U134 ( .A0(\b<4> ), .A1(n72), .B0(N17), .B1(n238), .Y(n71) );
  OAI2BB1X1 U135 ( .A0N(n241), .A1N(\a<4> ), .B0(n233), .Y(n72) );
  NAND2X1 U136 ( .A(n73), .B(n74), .Y(\Result<3> ) );
  AOI22X1 U137 ( .A0(N49), .A1(n229), .B0(\a<3> ), .B1(n232), .Y(n73) );
  AOI22X1 U138 ( .A0(\b<3> ), .A1(n75), .B0(N16), .B1(n238), .Y(n74) );
  OAI2BB1X1 U139 ( .A0N(n241), .A1N(\a<3> ), .B0(n233), .Y(n75) );
  NAND2X1 U140 ( .A(n85), .B(n86), .Y(\Result<6> ) );
  AOI22X1 U141 ( .A0(N52), .A1(n228), .B0(\a<6> ), .B1(n232), .Y(n85) );
  AOI22X1 U142 ( .A0(\b<6> ), .A1(n87), .B0(N19), .B1(n238), .Y(n86) );
  OAI2BB1X1 U143 ( .A0N(n241), .A1N(\a<6> ), .B0(n235), .Y(n87) );
  NAND2X1 U144 ( .A(n67), .B(n68), .Y(\Result<5> ) );
  AOI22X1 U145 ( .A0(N51), .A1(n229), .B0(\a<5> ), .B1(n232), .Y(n67) );
  AOI22X1 U146 ( .A0(\b<5> ), .A1(n69), .B0(N18), .B1(n238), .Y(n68) );
  OAI2BB1X1 U147 ( .A0N(n241), .A1N(\a<5> ), .B0(n235), .Y(n69) );
  OAI2BB1X1 U148 ( .A0N(n240), .A1N(\a<31> ), .B0(n235), .Y(n117) );
  AND2X2 U149 ( .A(\ALUControl<0> ), .B(n240), .Y(n226) );
  NAND2X1 U150 ( .A(n12), .B(n13), .Y(\Result<1> ) );
  AOI22X1 U151 ( .A0(N47), .A1(n228), .B0(\a<1> ), .B1(n232), .Y(n12) );
  AOI22X1 U152 ( .A0(\b<1> ), .A1(n14), .B0(N14), .B1(n238), .Y(n13) );
  OAI2BB1X1 U153 ( .A0N(n241), .A1N(\a<1> ), .B0(n236), .Y(n14) );
  NOR2BX1 U154 ( .AN(\ALUControl<0> ), .B(n240), .Y(n17) );
  NAND2X1 U155 ( .A(n48), .B(n49), .Y(\Result<0> ) );
  AOI22X1 U156 ( .A0(N46), .A1(n229), .B0(\a<0> ), .B1(n226), .Y(n48) );
  AOI22X1 U157 ( .A0(\b<0> ), .A1(n50), .B0(N13), .B1(n239), .Y(n49) );
  XOR2X1 U158 ( .A(\b<31> ), .B(\a<31> ), .Y(n114) );
  OAI2BB1X1 U159 ( .A0N(n241), .A1N(\a<0> ), .B0(n233), .Y(n50) );
  NOR2X1 U160 ( .A(n6), .B(n7), .Y(N173) );
  OR4X2 U161 ( .A(n8), .B(n9), .C(n10), .D(n11), .Y(n7) );
  NOR3X1 U162 ( .A(n112), .B(n240), .C(n113), .Y(\ALUFlags<0> ) );
  XOR2X1 U163 ( .A(\ALUControl<0> ), .B(n114), .Y(n113) );
  AND2X2 U164 ( .A(N45), .B(n239), .Y(\ALUFlags<1> ) );
  BUFX3 U165 ( .A(\Result<31> ), .Y(\ALUFlags<3> ) );
  NAND2X1 U166 ( .A(n115), .B(n116), .Y(\Result<31> ) );
endmodule


module datapath ( clk, reset, .Adr({\Adr<31> , \Adr<30> , \Adr<29> , \Adr<28> , 
        \Adr<27> , \Adr<26> , \Adr<25> , \Adr<24> , \Adr<23> , \Adr<22> , 
        \Adr<21> , \Adr<20> , \Adr<19> , \Adr<18> , \Adr<17> , \Adr<16> , 
        \Adr<15> , \Adr<14> , \Adr<13> , \Adr<12> , \Adr<11> , \Adr<10> , 
        \Adr<9> , \Adr<8> , \Adr<7> , \Adr<6> , \Adr<5> , \Adr<4> , \Adr<3> , 
        \Adr<2> , \Adr<1> , \Adr<0> }), .WriteData({\WriteData<31> , 
        \WriteData<30> , \WriteData<29> , \WriteData<28> , \WriteData<27> , 
        \WriteData<26> , \WriteData<25> , \WriteData<24> , \WriteData<23> , 
        \WriteData<22> , \WriteData<21> , \WriteData<20> , \WriteData<19> , 
        \WriteData<18> , \WriteData<17> , \WriteData<16> , \WriteData<15> , 
        \WriteData<14> , \WriteData<13> , \WriteData<12> , \WriteData<11> , 
        \WriteData<10> , \WriteData<9> , \WriteData<8> , \WriteData<7> , 
        \WriteData<6> , \WriteData<5> , \WriteData<4> , \WriteData<3> , 
        \WriteData<2> , \WriteData<1> , \WriteData<0> }), .ReadData({
        \ReadData<31> , \ReadData<30> , \ReadData<29> , \ReadData<28> , 
        \ReadData<27> , \ReadData<26> , \ReadData<25> , \ReadData<24> , 
        \ReadData<23> , \ReadData<22> , \ReadData<21> , \ReadData<20> , 
        \ReadData<19> , \ReadData<18> , \ReadData<17> , \ReadData<16> , 
        \ReadData<15> , \ReadData<14> , \ReadData<13> , \ReadData<12> , 
        \ReadData<11> , \ReadData<10> , \ReadData<9> , \ReadData<8> , 
        \ReadData<7> , \ReadData<6> , \ReadData<5> , \ReadData<4> , 
        \ReadData<3> , \ReadData<2> , \ReadData<1> , \ReadData<0> }), .Instr({
        \Instr<31> , \Instr<30> , \Instr<29> , \Instr<28> , \Instr<27> , 
        \Instr<26> , \Instr<25> , \Instr<24> , \Instr<23> , \Instr<22> , 
        \Instr<21> , \Instr<20> , \Instr<19> , \Instr<18> , \Instr<17> , 
        \Instr<16> , \Instr<15> , \Instr<14> , \Instr<13> , \Instr<12> , 
        \Instr<11> , \Instr<10> , \Instr<9> , \Instr<8> , \Instr<7> , 
        \Instr<6> , \Instr<5> , \Instr<4> , \Instr<3> , \Instr<2> , \Instr<1> , 
        \Instr<0> }), .ALUFlags({\ALUFlags<3> , \ALUFlags<2> , \ALUFlags<1> , 
        \ALUFlags<0> }), PCWrite, RegWrite, IRWrite, AdrSrc, .RegSrc({
        \RegSrc<1> , \RegSrc<0> }), .ALUSrcA({\ALUSrcA<1> , \ALUSrcA<0> }), 
    .ALUSrcB({\ALUSrcB<1> , \ALUSrcB<0> }), .ResultSrc({\ResultSrc<1> , 
        \ResultSrc<0> }), .ImmSrc({\ImmSrc<1> , \ImmSrc<0> }), .ALUControl({
        \ALUControl<1> , \ALUControl<0> }) );
  input clk, reset, \ReadData<31> , \ReadData<30> , \ReadData<29> ,
         \ReadData<28> , \ReadData<27> , \ReadData<26> , \ReadData<25> ,
         \ReadData<24> , \ReadData<23> , \ReadData<22> , \ReadData<21> ,
         \ReadData<20> , \ReadData<19> , \ReadData<18> , \ReadData<17> ,
         \ReadData<16> , \ReadData<15> , \ReadData<14> , \ReadData<13> ,
         \ReadData<12> , \ReadData<11> , \ReadData<10> , \ReadData<9> ,
         \ReadData<8> , \ReadData<7> , \ReadData<6> , \ReadData<5> ,
         \ReadData<4> , \ReadData<3> , \ReadData<2> , \ReadData<1> ,
         \ReadData<0> , PCWrite, RegWrite, IRWrite, AdrSrc, \RegSrc<1> ,
         \RegSrc<0> , \ALUSrcA<1> , \ALUSrcA<0> , \ALUSrcB<1> , \ALUSrcB<0> ,
         \ResultSrc<1> , \ResultSrc<0> , \ImmSrc<1> , \ImmSrc<0> ,
         \ALUControl<1> , \ALUControl<0> ;
  output \Adr<31> , \Adr<30> , \Adr<29> , \Adr<28> , \Adr<27> , \Adr<26> ,
         \Adr<25> , \Adr<24> , \Adr<23> , \Adr<22> , \Adr<21> , \Adr<20> ,
         \Adr<19> , \Adr<18> , \Adr<17> , \Adr<16> , \Adr<15> , \Adr<14> ,
         \Adr<13> , \Adr<12> , \Adr<11> , \Adr<10> , \Adr<9> , \Adr<8> ,
         \Adr<7> , \Adr<6> , \Adr<5> , \Adr<4> , \Adr<3> , \Adr<2> , \Adr<1> ,
         \Adr<0> , \WriteData<31> , \WriteData<30> , \WriteData<29> ,
         \WriteData<28> , \WriteData<27> , \WriteData<26> , \WriteData<25> ,
         \WriteData<24> , \WriteData<23> , \WriteData<22> , \WriteData<21> ,
         \WriteData<20> , \WriteData<19> , \WriteData<18> , \WriteData<17> ,
         \WriteData<16> , \WriteData<15> , \WriteData<14> , \WriteData<13> ,
         \WriteData<12> , \WriteData<11> , \WriteData<10> , \WriteData<9> ,
         \WriteData<8> , \WriteData<7> , \WriteData<6> , \WriteData<5> ,
         \WriteData<4> , \WriteData<3> , \WriteData<2> , \WriteData<1> ,
         \WriteData<0> , \Instr<31> , \Instr<30> , \Instr<29> , \Instr<28> ,
         \Instr<27> , \Instr<26> , \Instr<25> , \Instr<24> , \Instr<23> ,
         \Instr<22> , \Instr<21> , \Instr<20> , \Instr<19> , \Instr<18> ,
         \Instr<17> , \Instr<16> , \Instr<15> , \Instr<14> , \Instr<13> ,
         \Instr<12> , \Instr<11> , \Instr<10> , \Instr<9> , \Instr<8> ,
         \Instr<7> , \Instr<6> , \Instr<5> , \Instr<4> , \Instr<3> ,
         \Instr<2> , \Instr<1> , \Instr<0> , \ALUFlags<3> , \ALUFlags<2> ,
         \ALUFlags<1> , \ALUFlags<0> ;
  wire   \PC<31> , \PC<30> , \PC<29> , \PC<28> , \PC<27> , \PC<26> , \PC<25> ,
         \PC<24> , \PC<23> , \PC<22> , \PC<21> , \PC<20> , \PC<19> , \PC<18> ,
         \PC<17> , \PC<16> , \PC<15> , \PC<14> , \PC<13> , \PC<12> , \PC<11> ,
         \PC<10> , \PC<9> , \PC<8> , \PC<7> , \PC<6> , \PC<5> , \PC<4> ,
         \PC<3> , \PC<2> , \PC<1> , \PC<0> , \Data<31> , \Data<30> ,
         \Data<29> , \Data<28> , \Data<27> , \Data<26> , \Data<25> ,
         \Data<24> , \Data<23> , \Data<22> , \Data<21> , \Data<20> ,
         \Data<19> , \Data<18> , \Data<17> , \Data<16> , \Data<15> ,
         \Data<14> , \Data<13> , \Data<12> , \Data<11> , \Data<10> , \Data<9> ,
         \Data<8> , \Data<7> , \Data<6> , \Data<5> , \Data<4> , \Data<3> ,
         \Data<2> , \Data<1> , \Data<0> , \RD1<31> , \RD1<30> , \RD1<29> ,
         \RD1<28> , \RD1<27> , \RD1<26> , \RD1<25> , \RD1<24> , \RD1<23> ,
         \RD1<22> , \RD1<21> , \RD1<20> , \RD1<19> , \RD1<18> , \RD1<17> ,
         \RD1<16> , \RD1<15> , \RD1<14> , \RD1<13> , \RD1<12> , \RD1<11> ,
         \RD1<10> , \RD1<9> , \RD1<8> , \RD1<7> , \RD1<6> , \RD1<5> , \RD1<4> ,
         \RD1<3> , \RD1<2> , \RD1<1> , \RD1<0> , \A<31> , \A<30> , \A<29> ,
         \A<28> , \A<27> , \A<26> , \A<25> , \A<24> , \A<23> , \A<22> ,
         \A<21> , \A<20> , \A<19> , \A<18> , \A<17> , \A<16> , \A<15> ,
         \A<14> , \A<13> , \A<12> , \A<11> , \A<10> , \A<9> , \A<8> , \A<7> ,
         \A<6> , \A<5> , \A<4> , \A<3> , \A<2> , \A<1> , \A<0> , \RD2<31> ,
         \RD2<30> , \RD2<29> , \RD2<28> , \RD2<27> , \RD2<26> , \RD2<25> ,
         \RD2<24> , \RD2<23> , \RD2<22> , \RD2<21> , \RD2<20> , \RD2<19> ,
         \RD2<18> , \RD2<17> , \RD2<16> , \RD2<15> , \RD2<14> , \RD2<13> ,
         \RD2<12> , \RD2<11> , \RD2<10> , \RD2<9> , \RD2<8> , \RD2<7> ,
         \RD2<6> , \RD2<5> , \RD2<4> , \RD2<3> , \RD2<2> , \RD2<1> , \RD2<0> ,
         \ALUResult<31> , \ALUResult<30> , \ALUResult<29> , \ALUResult<28> ,
         \ALUResult<27> , \ALUResult<26> , \ALUResult<25> , \ALUResult<24> ,
         \ALUResult<23> , \ALUResult<22> , \ALUResult<21> , \ALUResult<20> ,
         \ALUResult<19> , \ALUResult<18> , \ALUResult<17> , \ALUResult<16> ,
         \ALUResult<15> , \ALUResult<14> , \ALUResult<13> , \ALUResult<12> ,
         \ALUResult<11> , \ALUResult<10> , \ALUResult<9> , \ALUResult<8> ,
         \ALUResult<7> , \ALUResult<6> , \ALUResult<5> , \ALUResult<4> ,
         \ALUResult<3> , \ALUResult<2> , \ALUResult<1> , \ALUResult<0> ,
         \ALUOut<31> , \ALUOut<30> , \ALUOut<29> , \ALUOut<28> , \ALUOut<27> ,
         \ALUOut<26> , \ALUOut<25> , \ALUOut<24> , \ALUOut<23> , \ALUOut<22> ,
         \ALUOut<21> , \ALUOut<20> , \ALUOut<19> , \ALUOut<18> , \ALUOut<17> ,
         \ALUOut<16> , \ALUOut<15> , \ALUOut<14> , \ALUOut<13> , \ALUOut<12> ,
         \ALUOut<11> , \ALUOut<10> , \ALUOut<9> , \ALUOut<8> , \ALUOut<7> ,
         \ALUOut<6> , \ALUOut<5> , \ALUOut<4> , \ALUOut<3> , \ALUOut<2> ,
         \ALUOut<1> , \ALUOut<0> , \Result<31> , \Result<30> , \Result<29> ,
         \Result<28> , \Result<27> , \Result<26> , \Result<25> , \Result<24> ,
         \Result<23> , \Result<22> , \Result<21> , \Result<20> , \Result<19> ,
         \Result<18> , \Result<17> , \Result<16> , \Result<15> , \Result<14> ,
         \Result<13> , \Result<12> , \Result<11> , \Result<10> , \Result<9> ,
         \Result<8> , \Result<7> , \Result<6> , \Result<5> , \Result<4> ,
         \Result<3> , \Result<2> , \Result<1> , \Result<0> , \RA1<3> ,
         \RA1<2> , \RA1<1> , \RA1<0> , \RA2<3> , \RA2<2> , \RA2<1> , \RA2<0> ,
         \SrcA<31> , \SrcA<30> , \SrcA<29> , \SrcA<28> , \SrcA<27> ,
         \SrcA<26> , \SrcA<25> , \SrcA<24> , \SrcA<23> , \SrcA<22> ,
         \SrcA<21> , \SrcA<20> , \SrcA<19> , \SrcA<18> , \SrcA<17> ,
         \SrcA<16> , \SrcA<15> , \SrcA<14> , \SrcA<13> , \SrcA<12> ,
         \SrcA<11> , \SrcA<10> , \SrcA<9> , \SrcA<8> , \SrcA<7> , \SrcA<6> ,
         \SrcA<5> , \SrcA<4> , \SrcA<3> , \SrcA<2> , \SrcA<1> , \SrcA<0> ,
         \ExtImm<31> , \ExtImm<30> , \ExtImm<29> , \ExtImm<28> , \ExtImm<27> ,
         \ExtImm<26> , \ExtImm<25> , \ExtImm<24> , \ExtImm<23> , \ExtImm<22> ,
         \ExtImm<21> , \ExtImm<20> , \ExtImm<19> , \ExtImm<18> , \ExtImm<17> ,
         \ExtImm<16> , \ExtImm<15> , \ExtImm<14> , \ExtImm<13> , \ExtImm<12> ,
         \ExtImm<11> , \ExtImm<10> , \ExtImm<9> , \ExtImm<8> , \ExtImm<7> ,
         \ExtImm<6> , \ExtImm<5> , \ExtImm<4> , \ExtImm<3> , \ExtImm<2> ,
         \ExtImm<1> , \ExtImm<0> , \SrcB<31> , \SrcB<30> , \SrcB<29> ,
         \SrcB<28> , \SrcB<27> , \SrcB<26> , \SrcB<25> , \SrcB<24> ,
         \SrcB<23> , \SrcB<22> , \SrcB<21> , \SrcB<20> , \SrcB<19> ,
         \SrcB<18> , \SrcB<17> , \SrcB<16> , \SrcB<15> , \SrcB<14> ,
         \SrcB<13> , \SrcB<12> , \SrcB<11> , \SrcB<10> , \SrcB<9> , \SrcB<8> ,
         \SrcB<7> , \SrcB<6> , \SrcB<5> , \SrcB<4> , \SrcB<3> , \SrcB<2> ,
         \SrcB<1> , \SrcB<0> , n787, n788, n789, n790, n791, n792, n793, n794,
         n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805,
         n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816,
         n817, n818, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n724, n726, n728, n730,
         n732, n734, n736, n738, n740, n742, n744, n746, n748, n750, n752,
         n754, n756, n758, n760, n762, n764, n766, n768, n770, n772, n774,
         n776, n778, n780, n782, n784, n786;

  flopenr_WIDTH32_0 pcreg ( .clk(clk), .reset(reset), .en(n721), .d({
        \Result<31> , \Result<30> , \Result<29> , \Result<28> , \Result<27> , 
        \Result<26> , \Result<25> , \Result<24> , \Result<23> , \Result<22> , 
        \Result<21> , \Result<20> , \Result<19> , \Result<18> , \Result<17> , 
        \Result<16> , \Result<15> , \Result<14> , \Result<13> , \Result<12> , 
        \Result<11> , \Result<10> , \Result<9> , \Result<8> , \Result<7> , 
        \Result<6> , \Result<5> , \Result<4> , \Result<3> , \Result<2> , 
        \Result<1> , \Result<0> }), .q({\PC<31> , \PC<30> , \PC<29> , \PC<28> , 
        \PC<27> , \PC<26> , \PC<25> , \PC<24> , \PC<23> , \PC<22> , \PC<21> , 
        \PC<20> , \PC<19> , \PC<18> , \PC<17> , \PC<16> , \PC<15> , \PC<14> , 
        \PC<13> , \PC<12> , \PC<11> , \PC<10> , \PC<9> , \PC<8> , \PC<7> , 
        \PC<6> , \PC<5> , \PC<4> , \PC<3> , \PC<2> , \PC<1> , \PC<0> }) );
  flopenr_WIDTH32_1 instrreg ( .clk(clk), .reset(reset), .en(n719), .d({
        \ReadData<31> , \ReadData<30> , \ReadData<29> , \ReadData<28> , 
        \ReadData<27> , \ReadData<26> , \ReadData<25> , \ReadData<24> , 
        \ReadData<23> , \ReadData<22> , \ReadData<21> , \ReadData<20> , 
        \ReadData<19> , \ReadData<18> , \ReadData<17> , \ReadData<16> , 
        \ReadData<15> , \ReadData<14> , \ReadData<13> , \ReadData<12> , 
        \ReadData<11> , \ReadData<10> , \ReadData<9> , \ReadData<8> , 
        \ReadData<7> , \ReadData<6> , \ReadData<5> , \ReadData<4> , 
        \ReadData<3> , \ReadData<2> , \ReadData<1> , \ReadData<0> }), .q({
        \Instr<31> , \Instr<30> , \Instr<29> , \Instr<28> , \Instr<27> , 
        \Instr<26> , \Instr<25> , \Instr<24> , \Instr<23> , \Instr<22> , 
        \Instr<21> , \Instr<20> , \Instr<19> , \Instr<18> , \Instr<17> , 
        \Instr<16> , \Instr<15> , \Instr<14> , \Instr<13> , \Instr<12> , 
        \Instr<11> , \Instr<10> , \Instr<9> , \Instr<8> , \Instr<7> , 
        \Instr<6> , \Instr<5> , \Instr<4> , \Instr<3> , \Instr<2> , \Instr<1> , 
        \Instr<0> }) );
  flopr_WIDTH32_0 datareg ( .clk(clk), .reset(reset), .d({\ReadData<31> , 
        \ReadData<30> , \ReadData<29> , \ReadData<28> , \ReadData<27> , 
        \ReadData<26> , \ReadData<25> , \ReadData<24> , \ReadData<23> , 
        \ReadData<22> , \ReadData<21> , \ReadData<20> , \ReadData<19> , 
        \ReadData<18> , \ReadData<17> , \ReadData<16> , \ReadData<15> , 
        \ReadData<14> , \ReadData<13> , \ReadData<12> , \ReadData<11> , 
        \ReadData<10> , \ReadData<9> , \ReadData<8> , \ReadData<7> , 
        \ReadData<6> , \ReadData<5> , \ReadData<4> , \ReadData<3> , 
        \ReadData<2> , \ReadData<1> , \ReadData<0> }), .q({\Data<31> , 
        \Data<30> , \Data<29> , \Data<28> , \Data<27> , \Data<26> , \Data<25> , 
        \Data<24> , \Data<23> , \Data<22> , \Data<21> , \Data<20> , \Data<19> , 
        \Data<18> , \Data<17> , \Data<16> , \Data<15> , \Data<14> , \Data<13> , 
        \Data<12> , \Data<11> , \Data<10> , \Data<9> , \Data<8> , \Data<7> , 
        \Data<6> , \Data<5> , \Data<4> , \Data<3> , \Data<2> , \Data<1> , 
        \Data<0> }) );
  flopr_WIDTH32_3 rd1reg ( .clk(clk), .reset(reset), .d({\RD1<31> , \RD1<30> , 
        \RD1<29> , \RD1<28> , \RD1<27> , \RD1<26> , \RD1<25> , \RD1<24> , 
        \RD1<23> , \RD1<22> , \RD1<21> , \RD1<20> , \RD1<19> , \RD1<18> , 
        \RD1<17> , \RD1<16> , \RD1<15> , \RD1<14> , \RD1<13> , \RD1<12> , 
        \RD1<11> , \RD1<10> , \RD1<9> , \RD1<8> , \RD1<7> , \RD1<6> , \RD1<5> , 
        \RD1<4> , \RD1<3> , \RD1<2> , \RD1<1> , \RD1<0> }), .q({\A<31> , 
        \A<30> , \A<29> , \A<28> , \A<27> , \A<26> , \A<25> , \A<24> , \A<23> , 
        \A<22> , \A<21> , \A<20> , \A<19> , \A<18> , \A<17> , \A<16> , \A<15> , 
        \A<14> , \A<13> , \A<12> , \A<11> , \A<10> , \A<9> , \A<8> , \A<7> , 
        \A<6> , \A<5> , \A<4> , \A<3> , \A<2> , \A<1> , \A<0> }) );
  flopr_WIDTH32_2 rd2reg ( .clk(clk), .reset(reset), .d({\RD2<31> , \RD2<30> , 
        \RD2<29> , \RD2<28> , \RD2<27> , \RD2<26> , \RD2<25> , \RD2<24> , 
        \RD2<23> , \RD2<22> , \RD2<21> , \RD2<20> , \RD2<19> , \RD2<18> , 
        \RD2<17> , \RD2<16> , \RD2<15> , \RD2<14> , \RD2<13> , \RD2<12> , 
        \RD2<11> , \RD2<10> , \RD2<9> , \RD2<8> , \RD2<7> , \RD2<6> , \RD2<5> , 
        \RD2<4> , \RD2<3> , \RD2<2> , \RD2<1> , \RD2<0> }), .q({n787, n788, 
        n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, 
        n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, 
        n813, n814, n815, n816, n817, n818}) );
  flopr_WIDTH32_1 alureg ( .clk(clk), .reset(reset), .d({\ALUResult<31> , 
        \ALUResult<30> , \ALUResult<29> , \ALUResult<28> , \ALUResult<27> , 
        \ALUResult<26> , \ALUResult<25> , \ALUResult<24> , \ALUResult<23> , 
        \ALUResult<22> , \ALUResult<21> , \ALUResult<20> , \ALUResult<19> , 
        \ALUResult<18> , \ALUResult<17> , \ALUResult<16> , \ALUResult<15> , 
        \ALUResult<14> , \ALUResult<13> , \ALUResult<12> , \ALUResult<11> , 
        \ALUResult<10> , \ALUResult<9> , \ALUResult<8> , \ALUResult<7> , 
        \ALUResult<6> , \ALUResult<5> , \ALUResult<4> , \ALUResult<3> , 
        \ALUResult<2> , \ALUResult<1> , \ALUResult<0> }), .q({\ALUOut<31> , 
        \ALUOut<30> , \ALUOut<29> , \ALUOut<28> , \ALUOut<27> , \ALUOut<26> , 
        \ALUOut<25> , \ALUOut<24> , \ALUOut<23> , \ALUOut<22> , \ALUOut<21> , 
        \ALUOut<20> , \ALUOut<19> , \ALUOut<18> , \ALUOut<17> , \ALUOut<16> , 
        \ALUOut<15> , \ALUOut<14> , \ALUOut<13> , \ALUOut<12> , \ALUOut<11> , 
        \ALUOut<10> , \ALUOut<9> , \ALUOut<8> , \ALUOut<7> , \ALUOut<6> , 
        \ALUOut<5> , \ALUOut<4> , \ALUOut<3> , \ALUOut<2> , \ALUOut<1> , 
        \ALUOut<0> }) );
  mux2_WIDTH32 adrmux ( .d0({\PC<31> , \PC<30> , \PC<29> , \PC<28> , \PC<27> , 
        \PC<26> , \PC<25> , \PC<24> , \PC<23> , \PC<22> , \PC<21> , \PC<20> , 
        \PC<19> , \PC<18> , \PC<17> , \PC<16> , \PC<15> , \PC<14> , \PC<13> , 
        \PC<12> , \PC<11> , \PC<10> , \PC<9> , \PC<8> , \PC<7> , \PC<6> , 
        \PC<5> , \PC<4> , \PC<3> , \PC<2> , \PC<1> , \PC<0> }), .d1({
        \Result<31> , \Result<30> , \Result<29> , \Result<28> , \Result<27> , 
        \Result<26> , \Result<25> , \Result<24> , \Result<23> , \Result<22> , 
        \Result<21> , \Result<20> , \Result<19> , \Result<18> , \Result<17> , 
        \Result<16> , \Result<15> , \Result<14> , \Result<13> , \Result<12> , 
        \Result<11> , \Result<10> , \Result<9> , \Result<8> , \Result<7> , 
        \Result<6> , \Result<5> , \Result<4> , \Result<3> , \Result<2> , 
        \Result<1> , \Result<0> }), .s(n717), .y({\Adr<31> , \Adr<30> , 
        \Adr<29> , \Adr<28> , \Adr<27> , \Adr<26> , \Adr<25> , \Adr<24> , 
        \Adr<23> , \Adr<22> , \Adr<21> , \Adr<20> , \Adr<19> , \Adr<18> , 
        \Adr<17> , \Adr<16> , \Adr<15> , \Adr<14> , \Adr<13> , \Adr<12> , 
        \Adr<11> , \Adr<10> , \Adr<9> , \Adr<8> , \Adr<7> , \Adr<6> , \Adr<5> , 
        \Adr<4> , \Adr<3> , \Adr<2> , \Adr<1> , \Adr<0> }) );
  mux2_WIDTH4_0 ra1mux ( .d0({\Instr<19> , \Instr<18> , \Instr<17> , 
        \Instr<16> }), .d1({1'b1, 1'b1, 1'b1, 1'b1}), .s(\RegSrc<0> ), .y({
        \RA1<3> , \RA1<2> , \RA1<1> , \RA1<0> }) );
  mux2_WIDTH4_1 ra2mux ( .d0({\Instr<3> , \Instr<2> , \Instr<1> , \Instr<0> }), 
        .d1({\Instr<15> , \Instr<14> , \Instr<13> , \Instr<12> }), .s(
        \RegSrc<1> ), .y({\RA2<3> , \RA2<2> , \RA2<1> , \RA2<0> }) );
  mux3_WIDTH32_0 srcAmux ( .d0({\A<31> , \A<30> , \A<29> , \A<28> , \A<27> , 
        \A<26> , \A<25> , \A<24> , \A<23> , \A<22> , \A<21> , \A<20> , \A<19> , 
        \A<18> , \A<17> , \A<16> , \A<15> , \A<14> , \A<13> , \A<12> , \A<11> , 
        \A<10> , \A<9> , \A<8> , \A<7> , \A<6> , \A<5> , \A<4> , \A<3> , 
        \A<2> , \A<1> , \A<0> }), .d1({\PC<31> , \PC<30> , \PC<29> , \PC<28> , 
        \PC<27> , \PC<26> , \PC<25> , \PC<24> , \PC<23> , \PC<22> , \PC<21> , 
        \PC<20> , \PC<19> , \PC<18> , \PC<17> , \PC<16> , \PC<15> , \PC<14> , 
        \PC<13> , \PC<12> , \PC<11> , \PC<10> , \PC<9> , \PC<8> , \PC<7> , 
        \PC<6> , \PC<5> , \PC<4> , \PC<3> , \PC<2> , \PC<1> , \PC<0> }), .d2({
        \ALUOut<31> , \ALUOut<30> , \ALUOut<29> , \ALUOut<28> , \ALUOut<27> , 
        \ALUOut<26> , \ALUOut<25> , \ALUOut<24> , \ALUOut<23> , \ALUOut<22> , 
        \ALUOut<21> , \ALUOut<20> , \ALUOut<19> , \ALUOut<18> , \ALUOut<17> , 
        \ALUOut<16> , \ALUOut<15> , \ALUOut<14> , \ALUOut<13> , \ALUOut<12> , 
        \ALUOut<11> , \ALUOut<10> , \ALUOut<9> , \ALUOut<8> , \ALUOut<7> , 
        \ALUOut<6> , \ALUOut<5> , \ALUOut<4> , \ALUOut<3> , \ALUOut<2> , 
        \ALUOut<1> , \ALUOut<0> }), .s({n715, n713}), .y({\SrcA<31> , 
        \SrcA<30> , \SrcA<29> , \SrcA<28> , \SrcA<27> , \SrcA<26> , \SrcA<25> , 
        \SrcA<24> , \SrcA<23> , \SrcA<22> , \SrcA<21> , \SrcA<20> , \SrcA<19> , 
        \SrcA<18> , \SrcA<17> , \SrcA<16> , \SrcA<15> , \SrcA<14> , \SrcA<13> , 
        \SrcA<12> , \SrcA<11> , \SrcA<10> , \SrcA<9> , \SrcA<8> , \SrcA<7> , 
        \SrcA<6> , \SrcA<5> , \SrcA<4> , \SrcA<3> , \SrcA<2> , \SrcA<1> , 
        \SrcA<0> }) );
  mux3_WIDTH32_2 srcBmux ( .d0({\WriteData<31> , \WriteData<30> , 
        \WriteData<29> , \WriteData<28> , \WriteData<27> , \WriteData<26> , 
        \WriteData<25> , \WriteData<24> , \WriteData<23> , \WriteData<22> , 
        \WriteData<21> , \WriteData<20> , \WriteData<19> , \WriteData<18> , 
        \WriteData<17> , \WriteData<16> , \WriteData<15> , \WriteData<14> , 
        \WriteData<13> , \WriteData<12> , \WriteData<11> , \WriteData<10> , 
        \WriteData<9> , \WriteData<8> , \WriteData<7> , \WriteData<6> , 
        \WriteData<5> , \WriteData<4> , \WriteData<3> , \WriteData<2> , 
        \WriteData<1> , \WriteData<0> }), .d1({\ExtImm<31> , \ExtImm<30> , 
        \ExtImm<29> , \ExtImm<28> , \ExtImm<27> , \ExtImm<26> , \ExtImm<25> , 
        \ExtImm<24> , \ExtImm<23> , \ExtImm<22> , \ExtImm<21> , \ExtImm<20> , 
        \ExtImm<19> , \ExtImm<18> , \ExtImm<17> , \ExtImm<16> , \ExtImm<15> , 
        \ExtImm<14> , \ExtImm<13> , \ExtImm<12> , \ExtImm<11> , \ExtImm<10> , 
        \ExtImm<9> , \ExtImm<8> , \ExtImm<7> , \ExtImm<6> , \ExtImm<5> , 
        \ExtImm<4> , \ExtImm<3> , \ExtImm<2> , \ExtImm<1> , \ExtImm<0> }), 
        .d2({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0}), .s({n711, 
        \ALUSrcB<0> }), .y({\SrcB<31> , \SrcB<30> , \SrcB<29> , \SrcB<28> , 
        \SrcB<27> , \SrcB<26> , \SrcB<25> , \SrcB<24> , \SrcB<23> , \SrcB<22> , 
        \SrcB<21> , \SrcB<20> , \SrcB<19> , \SrcB<18> , \SrcB<17> , \SrcB<16> , 
        \SrcB<15> , \SrcB<14> , \SrcB<13> , \SrcB<12> , \SrcB<11> , \SrcB<10> , 
        \SrcB<9> , \SrcB<8> , \SrcB<7> , \SrcB<6> , \SrcB<5> , \SrcB<4> , 
        \SrcB<3> , \SrcB<2> , \SrcB<1> , \SrcB<0> }) );
  mux3_WIDTH32_1 alumux ( .d0({\ALUOut<31> , \ALUOut<30> , \ALUOut<29> , 
        \ALUOut<28> , \ALUOut<27> , \ALUOut<26> , \ALUOut<25> , \ALUOut<24> , 
        \ALUOut<23> , \ALUOut<22> , \ALUOut<21> , \ALUOut<20> , \ALUOut<19> , 
        \ALUOut<18> , \ALUOut<17> , \ALUOut<16> , \ALUOut<15> , \ALUOut<14> , 
        \ALUOut<13> , \ALUOut<12> , \ALUOut<11> , \ALUOut<10> , \ALUOut<9> , 
        \ALUOut<8> , \ALUOut<7> , \ALUOut<6> , \ALUOut<5> , \ALUOut<4> , 
        \ALUOut<3> , \ALUOut<2> , \ALUOut<1> , \ALUOut<0> }), .d1({\Data<31> , 
        \Data<30> , \Data<29> , \Data<28> , \Data<27> , \Data<26> , \Data<25> , 
        \Data<24> , \Data<23> , \Data<22> , \Data<21> , \Data<20> , \Data<19> , 
        \Data<18> , \Data<17> , \Data<16> , \Data<15> , \Data<14> , \Data<13> , 
        \Data<12> , \Data<11> , \Data<10> , \Data<9> , \Data<8> , \Data<7> , 
        \Data<6> , \Data<5> , \Data<4> , \Data<3> , \Data<2> , \Data<1> , 
        \Data<0> }), .d2({\ALUResult<31> , \ALUResult<30> , \ALUResult<29> , 
        \ALUResult<28> , \ALUResult<27> , \ALUResult<26> , \ALUResult<25> , 
        \ALUResult<24> , \ALUResult<23> , \ALUResult<22> , \ALUResult<21> , 
        \ALUResult<20> , \ALUResult<19> , \ALUResult<18> , \ALUResult<17> , 
        \ALUResult<16> , \ALUResult<15> , \ALUResult<14> , \ALUResult<13> , 
        \ALUResult<12> , \ALUResult<11> , \ALUResult<10> , \ALUResult<9> , 
        \ALUResult<8> , \ALUResult<7> , \ALUResult<6> , \ALUResult<5> , 
        \ALUResult<4> , \ALUResult<3> , \ALUResult<2> , \ALUResult<1> , 
        \ALUResult<0> }), .s({n709, \ResultSrc<0> }), .y({\Result<31> , 
        \Result<30> , \Result<29> , \Result<28> , \Result<27> , \Result<26> , 
        \Result<25> , \Result<24> , \Result<23> , \Result<22> , \Result<21> , 
        \Result<20> , \Result<19> , \Result<18> , \Result<17> , \Result<16> , 
        \Result<15> , \Result<14> , \Result<13> , \Result<12> , \Result<11> , 
        \Result<10> , \Result<9> , \Result<8> , \Result<7> , \Result<6> , 
        \Result<5> , \Result<4> , \Result<3> , \Result<2> , \Result<1> , 
        \Result<0> }) );
  regfile rf ( .clk(clk), .we3(RegWrite), .ra1({\RA1<3> , \RA1<2> , \RA1<1> , 
        \RA1<0> }), .ra2({\RA2<3> , \RA2<2> , \RA2<1> , \RA2<0> }), .wa3({
        \Instr<15> , \Instr<14> , \Instr<13> , \Instr<12> }), .wd3({
        \Result<31> , \Result<30> , \Result<29> , \Result<28> , \Result<27> , 
        \Result<26> , \Result<25> , \Result<24> , \Result<23> , \Result<22> , 
        \Result<21> , \Result<20> , \Result<19> , \Result<18> , \Result<17> , 
        \Result<16> , \Result<15> , \Result<14> , \Result<13> , \Result<12> , 
        \Result<11> , \Result<10> , \Result<9> , \Result<8> , \Result<7> , 
        \Result<6> , \Result<5> , \Result<4> , \Result<3> , \Result<2> , 
        \Result<1> , \Result<0> }), .r15({\Result<31> , \Result<30> , 
        \Result<29> , \Result<28> , \Result<27> , \Result<26> , \Result<25> , 
        \Result<24> , \Result<23> , \Result<22> , \Result<21> , \Result<20> , 
        \Result<19> , \Result<18> , \Result<17> , \Result<16> , \Result<15> , 
        \Result<14> , \Result<13> , \Result<12> , \Result<11> , \Result<10> , 
        \Result<9> , \Result<8> , \Result<7> , \Result<6> , \Result<5> , 
        \Result<4> , \Result<3> , \Result<2> , \Result<1> , \Result<0> }), 
        .rd1({\RD1<31> , \RD1<30> , \RD1<29> , \RD1<28> , \RD1<27> , \RD1<26> , 
        \RD1<25> , \RD1<24> , \RD1<23> , \RD1<22> , \RD1<21> , \RD1<20> , 
        \RD1<19> , \RD1<18> , \RD1<17> , \RD1<16> , \RD1<15> , \RD1<14> , 
        \RD1<13> , \RD1<12> , \RD1<11> , \RD1<10> , \RD1<9> , \RD1<8> , 
        \RD1<7> , \RD1<6> , \RD1<5> , \RD1<4> , \RD1<3> , \RD1<2> , \RD1<1> , 
        \RD1<0> }), .rd2({\RD2<31> , \RD2<30> , \RD2<29> , \RD2<28> , 
        \RD2<27> , \RD2<26> , \RD2<25> , \RD2<24> , \RD2<23> , \RD2<22> , 
        \RD2<21> , \RD2<20> , \RD2<19> , \RD2<18> , \RD2<17> , \RD2<16> , 
        \RD2<15> , \RD2<14> , \RD2<13> , \RD2<12> , \RD2<11> , \RD2<10> , 
        \RD2<9> , \RD2<8> , \RD2<7> , \RD2<6> , \RD2<5> , \RD2<4> , \RD2<3> , 
        \RD2<2> , \RD2<1> , \RD2<0> }) );
  extend ext ( .Instr({\Instr<23> , \Instr<22> , \Instr<21> , \Instr<20> , 
        \Instr<19> , \Instr<18> , \Instr<17> , \Instr<16> , \Instr<15> , 
        \Instr<14> , \Instr<13> , \Instr<12> , \Instr<11> , \Instr<10> , 
        \Instr<9> , \Instr<8> , \Instr<7> , \Instr<6> , \Instr<5> , \Instr<4> , 
        \Instr<3> , \Instr<2> , \Instr<1> , \Instr<0> }), .ImmSrc({\ImmSrc<1> , 
        \ImmSrc<0> }), .ExtImm({\ExtImm<31> , \ExtImm<30> , \ExtImm<29> , 
        \ExtImm<28> , \ExtImm<27> , \ExtImm<26> , \ExtImm<25> , \ExtImm<24> , 
        \ExtImm<23> , \ExtImm<22> , \ExtImm<21> , \ExtImm<20> , \ExtImm<19> , 
        \ExtImm<18> , \ExtImm<17> , \ExtImm<16> , \ExtImm<15> , \ExtImm<14> , 
        \ExtImm<13> , \ExtImm<12> , \ExtImm<11> , \ExtImm<10> , \ExtImm<9> , 
        \ExtImm<8> , \ExtImm<7> , \ExtImm<6> , \ExtImm<5> , \ExtImm<4> , 
        \ExtImm<3> , \ExtImm<2> , \ExtImm<1> , \ExtImm<0> }) );
  alu alu ( .a({\SrcA<31> , \SrcA<30> , \SrcA<29> , \SrcA<28> , \SrcA<27> , 
        \SrcA<26> , \SrcA<25> , \SrcA<24> , \SrcA<23> , \SrcA<22> , \SrcA<21> , 
        \SrcA<20> , \SrcA<19> , \SrcA<18> , \SrcA<17> , \SrcA<16> , \SrcA<15> , 
        \SrcA<14> , \SrcA<13> , \SrcA<12> , \SrcA<11> , \SrcA<10> , \SrcA<9> , 
        \SrcA<8> , \SrcA<7> , \SrcA<6> , \SrcA<5> , \SrcA<4> , \SrcA<3> , 
        \SrcA<2> , \SrcA<1> , \SrcA<0> }), .b({\SrcB<31> , \SrcB<30> , 
        \SrcB<29> , \SrcB<28> , \SrcB<27> , \SrcB<26> , \SrcB<25> , \SrcB<24> , 
        \SrcB<23> , \SrcB<22> , \SrcB<21> , \SrcB<20> , \SrcB<19> , \SrcB<18> , 
        \SrcB<17> , \SrcB<16> , \SrcB<15> , \SrcB<14> , \SrcB<13> , \SrcB<12> , 
        \SrcB<11> , \SrcB<10> , \SrcB<9> , \SrcB<8> , \SrcB<7> , \SrcB<6> , 
        \SrcB<5> , \SrcB<4> , \SrcB<3> , \SrcB<2> , \SrcB<1> , \SrcB<0> }), 
        .ALUControl({n707, \ALUControl<0> }), .Result({\ALUResult<31> , 
        \ALUResult<30> , \ALUResult<29> , \ALUResult<28> , \ALUResult<27> , 
        \ALUResult<26> , \ALUResult<25> , \ALUResult<24> , \ALUResult<23> , 
        \ALUResult<22> , \ALUResult<21> , \ALUResult<20> , \ALUResult<19> , 
        \ALUResult<18> , \ALUResult<17> , \ALUResult<16> , \ALUResult<15> , 
        \ALUResult<14> , \ALUResult<13> , \ALUResult<12> , \ALUResult<11> , 
        \ALUResult<10> , \ALUResult<9> , \ALUResult<8> , \ALUResult<7> , 
        \ALUResult<6> , \ALUResult<5> , \ALUResult<4> , \ALUResult<3> , 
        \ALUResult<2> , \ALUResult<1> , \ALUResult<0> }), .ALUFlags({
        \ALUFlags<3> , \ALUFlags<2> , \ALUFlags<1> , \ALUFlags<0> }) );
  INVX1 U3 ( .A(n712), .Y(n711) );
  INVX1 U4 ( .A(\ALUSrcB<1> ), .Y(n712) );
  INVX1 U5 ( .A(n714), .Y(n713) );
  INVX1 U6 ( .A(\ALUSrcA<0> ), .Y(n714) );
  INVX1 U7 ( .A(n716), .Y(n715) );
  INVX1 U8 ( .A(\ALUSrcA<1> ), .Y(n716) );
  INVX1 U9 ( .A(n710), .Y(n709) );
  INVX1 U10 ( .A(\ResultSrc<1> ), .Y(n710) );
  INVX1 U11 ( .A(n720), .Y(n719) );
  INVX1 U12 ( .A(IRWrite), .Y(n720) );
  INVX1 U13 ( .A(n708), .Y(n707) );
  INVX1 U14 ( .A(\ALUControl<1> ), .Y(n708) );
  INVX1 U15 ( .A(n718), .Y(n717) );
  INVX1 U16 ( .A(AdrSrc), .Y(n718) );
  INVX1 U17 ( .A(n722), .Y(n721) );
  INVX1 U18 ( .A(PCWrite), .Y(n722) );
  INVX1 U19 ( .A(n724), .Y(\WriteData<0> ) );
  INVX1 U20 ( .A(n818), .Y(n724) );
  INVX1 U21 ( .A(n726), .Y(\WriteData<1> ) );
  INVX1 U22 ( .A(n817), .Y(n726) );
  INVX1 U23 ( .A(n728), .Y(\WriteData<2> ) );
  INVX1 U24 ( .A(n816), .Y(n728) );
  INVX1 U25 ( .A(n730), .Y(\WriteData<3> ) );
  INVX1 U26 ( .A(n815), .Y(n730) );
  INVX1 U27 ( .A(n732), .Y(\WriteData<4> ) );
  INVX1 U28 ( .A(n814), .Y(n732) );
  INVX1 U29 ( .A(n734), .Y(\WriteData<5> ) );
  INVX1 U30 ( .A(n813), .Y(n734) );
  INVX1 U31 ( .A(n736), .Y(\WriteData<6> ) );
  INVX1 U32 ( .A(n812), .Y(n736) );
  INVX1 U33 ( .A(n738), .Y(\WriteData<7> ) );
  INVX1 U34 ( .A(n811), .Y(n738) );
  INVX1 U35 ( .A(n740), .Y(\WriteData<8> ) );
  INVX1 U36 ( .A(n810), .Y(n740) );
  INVX1 U37 ( .A(n744), .Y(\WriteData<10> ) );
  INVX1 U38 ( .A(n808), .Y(n744) );
  INVX1 U39 ( .A(n746), .Y(\WriteData<11> ) );
  INVX1 U40 ( .A(n807), .Y(n746) );
  INVX1 U41 ( .A(n742), .Y(\WriteData<9> ) );
  INVX1 U42 ( .A(n809), .Y(n742) );
  INVX1 U43 ( .A(n748), .Y(\WriteData<12> ) );
  INVX1 U44 ( .A(n806), .Y(n748) );
  INVX1 U45 ( .A(n750), .Y(\WriteData<13> ) );
  INVX1 U46 ( .A(n805), .Y(n750) );
  INVX1 U47 ( .A(n752), .Y(\WriteData<14> ) );
  INVX1 U48 ( .A(n804), .Y(n752) );
  INVX1 U49 ( .A(n754), .Y(\WriteData<15> ) );
  INVX1 U50 ( .A(n803), .Y(n754) );
  INVX1 U51 ( .A(n756), .Y(\WriteData<16> ) );
  INVX1 U52 ( .A(n802), .Y(n756) );
  INVX1 U53 ( .A(n758), .Y(\WriteData<17> ) );
  INVX1 U54 ( .A(n801), .Y(n758) );
  INVX1 U55 ( .A(n760), .Y(\WriteData<18> ) );
  INVX1 U56 ( .A(n800), .Y(n760) );
  INVX1 U57 ( .A(n762), .Y(\WriteData<19> ) );
  INVX1 U58 ( .A(n799), .Y(n762) );
  INVX1 U59 ( .A(n764), .Y(\WriteData<20> ) );
  INVX1 U60 ( .A(n798), .Y(n764) );
  INVX1 U61 ( .A(n766), .Y(\WriteData<21> ) );
  INVX1 U62 ( .A(n797), .Y(n766) );
  INVX1 U63 ( .A(n768), .Y(\WriteData<22> ) );
  INVX1 U64 ( .A(n796), .Y(n768) );
  INVX1 U65 ( .A(n770), .Y(\WriteData<23> ) );
  INVX1 U66 ( .A(n795), .Y(n770) );
  INVX1 U67 ( .A(n772), .Y(\WriteData<24> ) );
  INVX1 U68 ( .A(n794), .Y(n772) );
  INVX1 U69 ( .A(n774), .Y(\WriteData<25> ) );
  INVX1 U70 ( .A(n793), .Y(n774) );
  INVX1 U71 ( .A(n776), .Y(\WriteData<26> ) );
  INVX1 U72 ( .A(n792), .Y(n776) );
  INVX1 U73 ( .A(n778), .Y(\WriteData<27> ) );
  INVX1 U74 ( .A(n791), .Y(n778) );
  INVX1 U75 ( .A(n780), .Y(\WriteData<28> ) );
  INVX1 U76 ( .A(n790), .Y(n780) );
  INVX1 U77 ( .A(n782), .Y(\WriteData<29> ) );
  INVX1 U78 ( .A(n789), .Y(n782) );
  INVX1 U79 ( .A(n784), .Y(\WriteData<30> ) );
  INVX1 U80 ( .A(n788), .Y(n784) );
  INVX1 U81 ( .A(n786), .Y(\WriteData<31> ) );
  INVX1 U82 ( .A(n787), .Y(n786) );
endmodule


module arm ( clk, reset, MemWrite, .Adr({\Adr<31> , \Adr<30> , \Adr<29> , 
        \Adr<28> , \Adr<27> , \Adr<26> , \Adr<25> , \Adr<24> , \Adr<23> , 
        \Adr<22> , \Adr<21> , \Adr<20> , \Adr<19> , \Adr<18> , \Adr<17> , 
        \Adr<16> , \Adr<15> , \Adr<14> , \Adr<13> , \Adr<12> , \Adr<11> , 
        \Adr<10> , \Adr<9> , \Adr<8> , \Adr<7> , \Adr<6> , \Adr<5> , \Adr<4> , 
        \Adr<3> , \Adr<2> , \Adr<1> , \Adr<0> }), .WriteData({\WriteData<31> , 
        \WriteData<30> , \WriteData<29> , \WriteData<28> , \WriteData<27> , 
        \WriteData<26> , \WriteData<25> , \WriteData<24> , \WriteData<23> , 
        \WriteData<22> , \WriteData<21> , \WriteData<20> , \WriteData<19> , 
        \WriteData<18> , \WriteData<17> , \WriteData<16> , \WriteData<15> , 
        \WriteData<14> , \WriteData<13> , \WriteData<12> , \WriteData<11> , 
        \WriteData<10> , \WriteData<9> , \WriteData<8> , \WriteData<7> , 
        \WriteData<6> , \WriteData<5> , \WriteData<4> , \WriteData<3> , 
        \WriteData<2> , \WriteData<1> , \WriteData<0> }), .ReadData({
        \ReadData<31> , \ReadData<30> , \ReadData<29> , \ReadData<28> , 
        \ReadData<27> , \ReadData<26> , \ReadData<25> , \ReadData<24> , 
        \ReadData<23> , \ReadData<22> , \ReadData<21> , \ReadData<20> , 
        \ReadData<19> , \ReadData<18> , \ReadData<17> , \ReadData<16> , 
        \ReadData<15> , \ReadData<14> , \ReadData<13> , \ReadData<12> , 
        \ReadData<11> , \ReadData<10> , \ReadData<9> , \ReadData<8> , 
        \ReadData<7> , \ReadData<6> , \ReadData<5> , \ReadData<4> , 
        \ReadData<3> , \ReadData<2> , \ReadData<1> , \ReadData<0> }) );
  input clk, reset, \ReadData<31> , \ReadData<30> , \ReadData<29> ,
         \ReadData<28> , \ReadData<27> , \ReadData<26> , \ReadData<25> ,
         \ReadData<24> , \ReadData<23> , \ReadData<22> , \ReadData<21> ,
         \ReadData<20> , \ReadData<19> , \ReadData<18> , \ReadData<17> ,
         \ReadData<16> , \ReadData<15> , \ReadData<14> , \ReadData<13> ,
         \ReadData<12> , \ReadData<11> , \ReadData<10> , \ReadData<9> ,
         \ReadData<8> , \ReadData<7> , \ReadData<6> , \ReadData<5> ,
         \ReadData<4> , \ReadData<3> , \ReadData<2> , \ReadData<1> ,
         \ReadData<0> ;
  output MemWrite, \Adr<31> , \Adr<30> , \Adr<29> , \Adr<28> , \Adr<27> ,
         \Adr<26> , \Adr<25> , \Adr<24> , \Adr<23> , \Adr<22> , \Adr<21> ,
         \Adr<20> , \Adr<19> , \Adr<18> , \Adr<17> , \Adr<16> , \Adr<15> ,
         \Adr<14> , \Adr<13> , \Adr<12> , \Adr<11> , \Adr<10> , \Adr<9> ,
         \Adr<8> , \Adr<7> , \Adr<6> , \Adr<5> , \Adr<4> , \Adr<3> , \Adr<2> ,
         \Adr<1> , \Adr<0> , \WriteData<31> , \WriteData<30> , \WriteData<29> ,
         \WriteData<28> , \WriteData<27> , \WriteData<26> , \WriteData<25> ,
         \WriteData<24> , \WriteData<23> , \WriteData<22> , \WriteData<21> ,
         \WriteData<20> , \WriteData<19> , \WriteData<18> , \WriteData<17> ,
         \WriteData<16> , \WriteData<15> , \WriteData<14> , \WriteData<13> ,
         \WriteData<12> , \WriteData<11> , \WriteData<10> , \WriteData<9> ,
         \WriteData<8> , \WriteData<7> , \WriteData<6> , \WriteData<5> ,
         \WriteData<4> , \WriteData<3> , \WriteData<2> , \WriteData<1> ,
         \WriteData<0> ;
  wire   \Instr<31> , \Instr<30> , \Instr<29> , \Instr<28> , \Instr<27> ,
         \Instr<26> , \Instr<25> , \Instr<24> , \Instr<23> , \Instr<22> ,
         \Instr<21> , \Instr<20> , \Instr<19> , \Instr<18> , \Instr<17> ,
         \Instr<16> , \Instr<15> , \Instr<14> , \Instr<13> , \Instr<12> ,
         \ALUFlags<3> , \ALUFlags<2> , \ALUFlags<1> , \ALUFlags<0> , PCWrite,
         RegWrite, IRWrite, AdrSrc, \RegSrc<1> , \RegSrc<0> , \ALUSrcA<1> ,
         \ALUSrcA<0> , \ALUSrcB<0> , \ResultSrc<1> , \ResultSrc<0> ,
         \ImmSrc<1> , \ImmSrc<0> , \ALUControl<1> , \ALUControl<0> , n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
         n784, n785, n786, n787, n788, n789, n790, n791, n792, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n698, n700, n702, n704, n706, n708, n710, n712, n714, n716,
         n718, n720, n722, n724, n726, n728, n730, n732, n734, n736, n738,
         n740, n742, n744, n746, n748, n750, n752, n754, n756, n758, n760;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12;

  controller c ( .clk(clk), .reset(reset), .Instr({\Instr<31> , \Instr<30> , 
        \Instr<29> , \Instr<28> , \Instr<27> , \Instr<26> , \Instr<25> , 
        \Instr<24> , \Instr<23> , \Instr<22> , \Instr<21> , \Instr<20> , 
        \Instr<19> , \Instr<18> , \Instr<17> , \Instr<16> , \Instr<15> , 
        \Instr<14> , \Instr<13> , \Instr<12> }), .ALUFlags({\ALUFlags<3> , 
        \ALUFlags<2> , \ALUFlags<1> , \ALUFlags<0> }), .PCWrite(PCWrite), 
        .MemWrite(MemWrite), .RegWrite(RegWrite), .IRWrite(IRWrite), .AdrSrc(
        AdrSrc), .RegSrc({\RegSrc<1> , \RegSrc<0> }), .ALUSrcA({\ALUSrcA<1> , 
        \ALUSrcA<0> }), .ALUSrcB({SYNOPSYS_UNCONNECTED__0, \ALUSrcB<0> }), 
        .ResultSrc({\ResultSrc<1> , \ResultSrc<0> }), .ImmSrc({\ImmSrc<1> , 
        \ImmSrc<0> }), .ALUControl({\ALUControl<1> , \ALUControl<0> }) );
  datapath dp ( .clk(clk), .reset(reset), .Adr({\Adr<31> , \Adr<30> , 
        \Adr<29> , \Adr<28> , \Adr<27> , \Adr<26> , \Adr<25> , \Adr<24> , 
        \Adr<23> , \Adr<22> , \Adr<21> , \Adr<20> , \Adr<19> , \Adr<18> , 
        \Adr<17> , \Adr<16> , \Adr<15> , \Adr<14> , \Adr<13> , \Adr<12> , 
        \Adr<11> , \Adr<10> , \Adr<9> , \Adr<8> , \Adr<7> , \Adr<6> , \Adr<5> , 
        \Adr<4> , \Adr<3> , \Adr<2> , \Adr<1> , \Adr<0> }), .WriteData({n761, 
        n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, 
        n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, 
        n786, n787, n788, n789, n790, n791, n792}), .ReadData({\ReadData<31> , 
        \ReadData<30> , \ReadData<29> , \ReadData<28> , \ReadData<27> , 
        \ReadData<26> , \ReadData<25> , \ReadData<24> , \ReadData<23> , 
        \ReadData<22> , \ReadData<21> , \ReadData<20> , \ReadData<19> , 
        \ReadData<18> , \ReadData<17> , \ReadData<16> , \ReadData<15> , 
        \ReadData<14> , \ReadData<13> , \ReadData<12> , \ReadData<11> , 
        \ReadData<10> , \ReadData<9> , \ReadData<8> , \ReadData<7> , 
        \ReadData<6> , \ReadData<5> , \ReadData<4> , \ReadData<3> , 
        \ReadData<2> , \ReadData<1> , \ReadData<0> }), .Instr({\Instr<31> , 
        \Instr<30> , \Instr<29> , \Instr<28> , \Instr<27> , \Instr<26> , 
        \Instr<25> , \Instr<24> , \Instr<23> , \Instr<22> , \Instr<21> , 
        \Instr<20> , \Instr<19> , \Instr<18> , \Instr<17> , \Instr<16> , 
        \Instr<15> , \Instr<14> , \Instr<13> , \Instr<12> , 
        SYNOPSYS_UNCONNECTED__1, SYNOPSYS_UNCONNECTED__2, 
        SYNOPSYS_UNCONNECTED__3, SYNOPSYS_UNCONNECTED__4, 
        SYNOPSYS_UNCONNECTED__5, SYNOPSYS_UNCONNECTED__6, 
        SYNOPSYS_UNCONNECTED__7, SYNOPSYS_UNCONNECTED__8, 
        SYNOPSYS_UNCONNECTED__9, SYNOPSYS_UNCONNECTED__10, 
        SYNOPSYS_UNCONNECTED__11, SYNOPSYS_UNCONNECTED__12}), .ALUFlags({
        \ALUFlags<3> , \ALUFlags<2> , \ALUFlags<1> , \ALUFlags<0> }), 
        .PCWrite(n695), .RegWrite(RegWrite), .IRWrite(n693), .AdrSrc(n691), 
        .RegSrc({\RegSrc<1> , \RegSrc<0> }), .ALUSrcA({n689, n687}), .ALUSrcB(
        {n687, \ALUSrcB<0> }), .ResultSrc({n685, \ResultSrc<0> }), .ImmSrc({
        \ImmSrc<1> , \ImmSrc<0> }), .ALUControl({n683, \ALUControl<0> }) );
  INVX1 U1 ( .A(n688), .Y(n687) );
  INVX1 U2 ( .A(\ALUSrcA<0> ), .Y(n688) );
  INVX1 U3 ( .A(n690), .Y(n689) );
  INVX1 U4 ( .A(\ALUSrcA<1> ), .Y(n690) );
  INVX1 U5 ( .A(n686), .Y(n685) );
  INVX1 U6 ( .A(\ResultSrc<1> ), .Y(n686) );
  INVX1 U7 ( .A(n692), .Y(n691) );
  INVX1 U8 ( .A(n694), .Y(n693) );
  INVX1 U9 ( .A(IRWrite), .Y(n694) );
  INVX1 U10 ( .A(n684), .Y(n683) );
  INVX1 U11 ( .A(\ALUControl<1> ), .Y(n684) );
  INVX1 U12 ( .A(AdrSrc), .Y(n692) );
  INVX1 U13 ( .A(n696), .Y(n695) );
  INVX1 U14 ( .A(PCWrite), .Y(n696) );
  INVX1 U15 ( .A(n698), .Y(\WriteData<0> ) );
  INVX1 U16 ( .A(n792), .Y(n698) );
  INVX1 U17 ( .A(n700), .Y(\WriteData<1> ) );
  INVX1 U18 ( .A(n791), .Y(n700) );
  INVX1 U19 ( .A(n702), .Y(\WriteData<2> ) );
  INVX1 U20 ( .A(n790), .Y(n702) );
  INVX1 U21 ( .A(n704), .Y(\WriteData<3> ) );
  INVX1 U22 ( .A(n789), .Y(n704) );
  INVX1 U23 ( .A(n706), .Y(\WriteData<4> ) );
  INVX1 U24 ( .A(n788), .Y(n706) );
  INVX1 U25 ( .A(n708), .Y(\WriteData<5> ) );
  INVX1 U26 ( .A(n787), .Y(n708) );
  INVX1 U27 ( .A(n710), .Y(\WriteData<6> ) );
  INVX1 U28 ( .A(n786), .Y(n710) );
  INVX1 U29 ( .A(n712), .Y(\WriteData<7> ) );
  INVX1 U30 ( .A(n785), .Y(n712) );
  INVX1 U31 ( .A(n714), .Y(\WriteData<8> ) );
  INVX1 U32 ( .A(n784), .Y(n714) );
  INVX1 U33 ( .A(n716), .Y(\WriteData<9> ) );
  INVX1 U34 ( .A(n783), .Y(n716) );
  INVX1 U35 ( .A(n718), .Y(\WriteData<10> ) );
  INVX1 U36 ( .A(n782), .Y(n718) );
  INVX1 U37 ( .A(n720), .Y(\WriteData<11> ) );
  INVX1 U38 ( .A(n781), .Y(n720) );
  INVX1 U39 ( .A(n722), .Y(\WriteData<12> ) );
  INVX1 U40 ( .A(n780), .Y(n722) );
  INVX1 U41 ( .A(n724), .Y(\WriteData<13> ) );
  INVX1 U42 ( .A(n779), .Y(n724) );
  INVX1 U43 ( .A(n726), .Y(\WriteData<14> ) );
  INVX1 U44 ( .A(n778), .Y(n726) );
  INVX1 U45 ( .A(n728), .Y(\WriteData<15> ) );
  INVX1 U46 ( .A(n777), .Y(n728) );
  INVX1 U47 ( .A(n730), .Y(\WriteData<16> ) );
  INVX1 U48 ( .A(n776), .Y(n730) );
  INVX1 U49 ( .A(n732), .Y(\WriteData<17> ) );
  INVX1 U50 ( .A(n775), .Y(n732) );
  INVX1 U51 ( .A(n734), .Y(\WriteData<18> ) );
  INVX1 U52 ( .A(n774), .Y(n734) );
  INVX1 U53 ( .A(n736), .Y(\WriteData<19> ) );
  INVX1 U54 ( .A(n773), .Y(n736) );
  INVX1 U55 ( .A(n738), .Y(\WriteData<20> ) );
  INVX1 U56 ( .A(n772), .Y(n738) );
  INVX1 U57 ( .A(n740), .Y(\WriteData<21> ) );
  INVX1 U58 ( .A(n771), .Y(n740) );
  INVX1 U59 ( .A(n742), .Y(\WriteData<22> ) );
  INVX1 U60 ( .A(n770), .Y(n742) );
  INVX1 U61 ( .A(n744), .Y(\WriteData<23> ) );
  INVX1 U62 ( .A(n769), .Y(n744) );
  INVX1 U63 ( .A(n746), .Y(\WriteData<24> ) );
  INVX1 U64 ( .A(n768), .Y(n746) );
  INVX1 U65 ( .A(n748), .Y(\WriteData<25> ) );
  INVX1 U66 ( .A(n767), .Y(n748) );
  INVX1 U67 ( .A(n750), .Y(\WriteData<26> ) );
  INVX1 U68 ( .A(n766), .Y(n750) );
  INVX1 U69 ( .A(n752), .Y(\WriteData<27> ) );
  INVX1 U70 ( .A(n765), .Y(n752) );
  INVX1 U71 ( .A(n754), .Y(\WriteData<28> ) );
  INVX1 U72 ( .A(n764), .Y(n754) );
  INVX1 U73 ( .A(n756), .Y(\WriteData<29> ) );
  INVX1 U74 ( .A(n763), .Y(n756) );
  INVX1 U75 ( .A(n758), .Y(\WriteData<30> ) );
  INVX1 U76 ( .A(n762), .Y(n758) );
  INVX1 U77 ( .A(n760), .Y(\WriteData<31> ) );
  INVX1 U78 ( .A(n761), .Y(n760) );
endmodule


module mem ( clk, we, .a({\a<31> , \a<30> , \a<29> , \a<28> , \a<27> , \a<26> , 
        \a<25> , \a<24> , \a<23> , \a<22> , \a<21> , \a<20> , \a<19> , \a<18> , 
        \a<17> , \a<16> , \a<15> , \a<14> , \a<13> , \a<12> , \a<11> , \a<10> , 
        \a<9> , \a<8> , \a<7> , \a<6> , \a<5> , \a<4> , \a<3> , \a<2> , \a<1> , 
        \a<0> }), .wd({\wd<31> , \wd<30> , \wd<29> , \wd<28> , \wd<27> , 
        \wd<26> , \wd<25> , \wd<24> , \wd<23> , \wd<22> , \wd<21> , \wd<20> , 
        \wd<19> , \wd<18> , \wd<17> , \wd<16> , \wd<15> , \wd<14> , \wd<13> , 
        \wd<12> , \wd<11> , \wd<10> , \wd<9> , \wd<8> , \wd<7> , \wd<6> , 
        \wd<5> , \wd<4> , \wd<3> , \wd<2> , \wd<1> , \wd<0> }), .rd({\rd<31> , 
        \rd<30> , \rd<29> , \rd<28> , \rd<27> , \rd<26> , \rd<25> , \rd<24> , 
        \rd<23> , \rd<22> , \rd<21> , \rd<20> , \rd<19> , \rd<18> , \rd<17> , 
        \rd<16> , \rd<15> , \rd<14> , \rd<13> , \rd<12> , \rd<11> , \rd<10> , 
        \rd<9> , \rd<8> , \rd<7> , \rd<6> , \rd<5> , \rd<4> , \rd<3> , \rd<2> , 
        \rd<1> , \rd<0> }) );
  input clk, we, \a<31> , \a<30> , \a<29> , \a<28> , \a<27> , \a<26> , \a<25> ,
         \a<24> , \a<23> , \a<22> , \a<21> , \a<20> , \a<19> , \a<18> ,
         \a<17> , \a<16> , \a<15> , \a<14> , \a<13> , \a<12> , \a<11> ,
         \a<10> , \a<9> , \a<8> , \a<7> , \a<6> , \a<5> , \a<4> , \a<3> ,
         \a<2> , \a<1> , \a<0> , \wd<31> , \wd<30> , \wd<29> , \wd<28> ,
         \wd<27> , \wd<26> , \wd<25> , \wd<24> , \wd<23> , \wd<22> , \wd<21> ,
         \wd<20> , \wd<19> , \wd<18> , \wd<17> , \wd<16> , \wd<15> , \wd<14> ,
         \wd<13> , \wd<12> , \wd<11> , \wd<10> , \wd<9> , \wd<8> , \wd<7> ,
         \wd<6> , \wd<5> , \wd<4> , \wd<3> , \wd<2> , \wd<1> , \wd<0> ;
  output \rd<31> , \rd<30> , \rd<29> , \rd<28> , \rd<27> , \rd<26> , \rd<25> ,
         \rd<24> , \rd<23> , \rd<22> , \rd<21> , \rd<20> , \rd<19> , \rd<18> ,
         \rd<17> , \rd<16> , \rd<15> , \rd<14> , \rd<13> , \rd<12> , \rd<11> ,
         \rd<10> , \rd<9> , \rd<8> , \rd<7> , \rd<6> , \rd<5> , \rd<4> ,
         \rd<3> , \rd<2> , \rd<1> , \rd<0> ;
  wire   N32, N33, N34, N35, N36, N37, \RAM<63><31> , \RAM<63><30> ,
         \RAM<63><29> , \RAM<63><28> , \RAM<63><27> , \RAM<63><26> ,
         \RAM<63><25> , \RAM<63><24> , \RAM<63><23> , \RAM<63><22> ,
         \RAM<63><21> , \RAM<63><20> , \RAM<63><19> , \RAM<63><18> ,
         \RAM<63><17> , \RAM<63><16> , \RAM<63><15> , \RAM<63><14> ,
         \RAM<63><13> , \RAM<63><12> , \RAM<63><11> , \RAM<63><10> ,
         \RAM<63><9> , \RAM<63><8> , \RAM<63><7> , \RAM<63><6> , \RAM<63><5> ,
         \RAM<63><4> , \RAM<63><3> , \RAM<63><2> , \RAM<63><1> , \RAM<63><0> ,
         \RAM<62><31> , \RAM<62><30> , \RAM<62><29> , \RAM<62><28> ,
         \RAM<62><27> , \RAM<62><26> , \RAM<62><25> , \RAM<62><24> ,
         \RAM<62><23> , \RAM<62><22> , \RAM<62><21> , \RAM<62><20> ,
         \RAM<62><19> , \RAM<62><18> , \RAM<62><17> , \RAM<62><16> ,
         \RAM<62><15> , \RAM<62><14> , \RAM<62><13> , \RAM<62><12> ,
         \RAM<62><11> , \RAM<62><10> , \RAM<62><9> , \RAM<62><8> ,
         \RAM<62><7> , \RAM<62><6> , \RAM<62><5> , \RAM<62><4> , \RAM<62><3> ,
         \RAM<62><2> , \RAM<62><1> , \RAM<62><0> , \RAM<61><31> ,
         \RAM<61><30> , \RAM<61><29> , \RAM<61><28> , \RAM<61><27> ,
         \RAM<61><26> , \RAM<61><25> , \RAM<61><24> , \RAM<61><23> ,
         \RAM<61><22> , \RAM<61><21> , \RAM<61><20> , \RAM<61><19> ,
         \RAM<61><18> , \RAM<61><17> , \RAM<61><16> , \RAM<61><15> ,
         \RAM<61><14> , \RAM<61><13> , \RAM<61><12> , \RAM<61><11> ,
         \RAM<61><10> , \RAM<61><9> , \RAM<61><8> , \RAM<61><7> , \RAM<61><6> ,
         \RAM<61><5> , \RAM<61><4> , \RAM<61><3> , \RAM<61><2> , \RAM<61><1> ,
         \RAM<61><0> , \RAM<60><31> , \RAM<60><30> , \RAM<60><29> ,
         \RAM<60><28> , \RAM<60><27> , \RAM<60><26> , \RAM<60><25> ,
         \RAM<60><24> , \RAM<60><23> , \RAM<60><22> , \RAM<60><21> ,
         \RAM<60><20> , \RAM<60><19> , \RAM<60><18> , \RAM<60><17> ,
         \RAM<60><16> , \RAM<60><15> , \RAM<60><14> , \RAM<60><13> ,
         \RAM<60><12> , \RAM<60><11> , \RAM<60><10> , \RAM<60><9> ,
         \RAM<60><8> , \RAM<60><7> , \RAM<60><6> , \RAM<60><5> , \RAM<60><4> ,
         \RAM<60><3> , \RAM<60><2> , \RAM<60><1> , \RAM<60><0> , \RAM<59><31> ,
         \RAM<59><30> , \RAM<59><29> , \RAM<59><28> , \RAM<59><27> ,
         \RAM<59><26> , \RAM<59><25> , \RAM<59><24> , \RAM<59><23> ,
         \RAM<59><22> , \RAM<59><21> , \RAM<59><20> , \RAM<59><19> ,
         \RAM<59><18> , \RAM<59><17> , \RAM<59><16> , \RAM<59><15> ,
         \RAM<59><14> , \RAM<59><13> , \RAM<59><12> , \RAM<59><11> ,
         \RAM<59><10> , \RAM<59><9> , \RAM<59><8> , \RAM<59><7> , \RAM<59><6> ,
         \RAM<59><5> , \RAM<59><4> , \RAM<59><3> , \RAM<59><2> , \RAM<59><1> ,
         \RAM<59><0> , \RAM<58><31> , \RAM<58><30> , \RAM<58><29> ,
         \RAM<58><28> , \RAM<58><27> , \RAM<58><26> , \RAM<58><25> ,
         \RAM<58><24> , \RAM<58><23> , \RAM<58><22> , \RAM<58><21> ,
         \RAM<58><20> , \RAM<58><19> , \RAM<58><18> , \RAM<58><17> ,
         \RAM<58><16> , \RAM<58><15> , \RAM<58><14> , \RAM<58><13> ,
         \RAM<58><12> , \RAM<58><11> , \RAM<58><10> , \RAM<58><9> ,
         \RAM<58><8> , \RAM<58><7> , \RAM<58><6> , \RAM<58><5> , \RAM<58><4> ,
         \RAM<58><3> , \RAM<58><2> , \RAM<58><1> , \RAM<58><0> , \RAM<57><31> ,
         \RAM<57><30> , \RAM<57><29> , \RAM<57><28> , \RAM<57><27> ,
         \RAM<57><26> , \RAM<57><25> , \RAM<57><24> , \RAM<57><23> ,
         \RAM<57><22> , \RAM<57><21> , \RAM<57><20> , \RAM<57><19> ,
         \RAM<57><18> , \RAM<57><17> , \RAM<57><16> , \RAM<57><15> ,
         \RAM<57><14> , \RAM<57><13> , \RAM<57><12> , \RAM<57><11> ,
         \RAM<57><10> , \RAM<57><9> , \RAM<57><8> , \RAM<57><7> , \RAM<57><6> ,
         \RAM<57><5> , \RAM<57><4> , \RAM<57><3> , \RAM<57><2> , \RAM<57><1> ,
         \RAM<57><0> , \RAM<56><31> , \RAM<56><30> , \RAM<56><29> ,
         \RAM<56><28> , \RAM<56><27> , \RAM<56><26> , \RAM<56><25> ,
         \RAM<56><24> , \RAM<56><23> , \RAM<56><22> , \RAM<56><21> ,
         \RAM<56><20> , \RAM<56><19> , \RAM<56><18> , \RAM<56><17> ,
         \RAM<56><16> , \RAM<56><15> , \RAM<56><14> , \RAM<56><13> ,
         \RAM<56><12> , \RAM<56><11> , \RAM<56><10> , \RAM<56><9> ,
         \RAM<56><8> , \RAM<56><7> , \RAM<56><6> , \RAM<56><5> , \RAM<56><4> ,
         \RAM<56><3> , \RAM<56><2> , \RAM<56><1> , \RAM<56><0> , \RAM<55><31> ,
         \RAM<55><30> , \RAM<55><29> , \RAM<55><28> , \RAM<55><27> ,
         \RAM<55><26> , \RAM<55><25> , \RAM<55><24> , \RAM<55><23> ,
         \RAM<55><22> , \RAM<55><21> , \RAM<55><20> , \RAM<55><19> ,
         \RAM<55><18> , \RAM<55><17> , \RAM<55><16> , \RAM<55><15> ,
         \RAM<55><14> , \RAM<55><13> , \RAM<55><12> , \RAM<55><11> ,
         \RAM<55><10> , \RAM<55><9> , \RAM<55><8> , \RAM<55><7> , \RAM<55><6> ,
         \RAM<55><5> , \RAM<55><4> , \RAM<55><3> , \RAM<55><2> , \RAM<55><1> ,
         \RAM<55><0> , \RAM<54><31> , \RAM<54><30> , \RAM<54><29> ,
         \RAM<54><28> , \RAM<54><27> , \RAM<54><26> , \RAM<54><25> ,
         \RAM<54><24> , \RAM<54><23> , \RAM<54><22> , \RAM<54><21> ,
         \RAM<54><20> , \RAM<54><19> , \RAM<54><18> , \RAM<54><17> ,
         \RAM<54><16> , \RAM<54><15> , \RAM<54><14> , \RAM<54><13> ,
         \RAM<54><12> , \RAM<54><11> , \RAM<54><10> , \RAM<54><9> ,
         \RAM<54><8> , \RAM<54><7> , \RAM<54><6> , \RAM<54><5> , \RAM<54><4> ,
         \RAM<54><3> , \RAM<54><2> , \RAM<54><1> , \RAM<54><0> , \RAM<53><31> ,
         \RAM<53><30> , \RAM<53><29> , \RAM<53><28> , \RAM<53><27> ,
         \RAM<53><26> , \RAM<53><25> , \RAM<53><24> , \RAM<53><23> ,
         \RAM<53><22> , \RAM<53><21> , \RAM<53><20> , \RAM<53><19> ,
         \RAM<53><18> , \RAM<53><17> , \RAM<53><16> , \RAM<53><15> ,
         \RAM<53><14> , \RAM<53><13> , \RAM<53><12> , \RAM<53><11> ,
         \RAM<53><10> , \RAM<53><9> , \RAM<53><8> , \RAM<53><7> , \RAM<53><6> ,
         \RAM<53><5> , \RAM<53><4> , \RAM<53><3> , \RAM<53><2> , \RAM<53><1> ,
         \RAM<53><0> , \RAM<52><31> , \RAM<52><30> , \RAM<52><29> ,
         \RAM<52><28> , \RAM<52><27> , \RAM<52><26> , \RAM<52><25> ,
         \RAM<52><24> , \RAM<52><23> , \RAM<52><22> , \RAM<52><21> ,
         \RAM<52><20> , \RAM<52><19> , \RAM<52><18> , \RAM<52><17> ,
         \RAM<52><16> , \RAM<52><15> , \RAM<52><14> , \RAM<52><13> ,
         \RAM<52><12> , \RAM<52><11> , \RAM<52><10> , \RAM<52><9> ,
         \RAM<52><8> , \RAM<52><7> , \RAM<52><6> , \RAM<52><5> , \RAM<52><4> ,
         \RAM<52><3> , \RAM<52><2> , \RAM<52><1> , \RAM<52><0> , \RAM<51><31> ,
         \RAM<51><30> , \RAM<51><29> , \RAM<51><28> , \RAM<51><27> ,
         \RAM<51><26> , \RAM<51><25> , \RAM<51><24> , \RAM<51><23> ,
         \RAM<51><22> , \RAM<51><21> , \RAM<51><20> , \RAM<51><19> ,
         \RAM<51><18> , \RAM<51><17> , \RAM<51><16> , \RAM<51><15> ,
         \RAM<51><14> , \RAM<51><13> , \RAM<51><12> , \RAM<51><11> ,
         \RAM<51><10> , \RAM<51><9> , \RAM<51><8> , \RAM<51><7> , \RAM<51><6> ,
         \RAM<51><5> , \RAM<51><4> , \RAM<51><3> , \RAM<51><2> , \RAM<51><1> ,
         \RAM<51><0> , \RAM<50><31> , \RAM<50><30> , \RAM<50><29> ,
         \RAM<50><28> , \RAM<50><27> , \RAM<50><26> , \RAM<50><25> ,
         \RAM<50><24> , \RAM<50><23> , \RAM<50><22> , \RAM<50><21> ,
         \RAM<50><20> , \RAM<50><19> , \RAM<50><18> , \RAM<50><17> ,
         \RAM<50><16> , \RAM<50><15> , \RAM<50><14> , \RAM<50><13> ,
         \RAM<50><12> , \RAM<50><11> , \RAM<50><10> , \RAM<50><9> ,
         \RAM<50><8> , \RAM<50><7> , \RAM<50><6> , \RAM<50><5> , \RAM<50><4> ,
         \RAM<50><3> , \RAM<50><2> , \RAM<50><1> , \RAM<50><0> , \RAM<49><31> ,
         \RAM<49><30> , \RAM<49><29> , \RAM<49><28> , \RAM<49><27> ,
         \RAM<49><26> , \RAM<49><25> , \RAM<49><24> , \RAM<49><23> ,
         \RAM<49><22> , \RAM<49><21> , \RAM<49><20> , \RAM<49><19> ,
         \RAM<49><18> , \RAM<49><17> , \RAM<49><16> , \RAM<49><15> ,
         \RAM<49><14> , \RAM<49><13> , \RAM<49><12> , \RAM<49><11> ,
         \RAM<49><10> , \RAM<49><9> , \RAM<49><8> , \RAM<49><7> , \RAM<49><6> ,
         \RAM<49><5> , \RAM<49><4> , \RAM<49><3> , \RAM<49><2> , \RAM<49><1> ,
         \RAM<49><0> , \RAM<48><31> , \RAM<48><30> , \RAM<48><29> ,
         \RAM<48><28> , \RAM<48><27> , \RAM<48><26> , \RAM<48><25> ,
         \RAM<48><24> , \RAM<48><23> , \RAM<48><22> , \RAM<48><21> ,
         \RAM<48><20> , \RAM<48><19> , \RAM<48><18> , \RAM<48><17> ,
         \RAM<48><16> , \RAM<48><15> , \RAM<48><14> , \RAM<48><13> ,
         \RAM<48><12> , \RAM<48><11> , \RAM<48><10> , \RAM<48><9> ,
         \RAM<48><8> , \RAM<48><7> , \RAM<48><6> , \RAM<48><5> , \RAM<48><4> ,
         \RAM<48><3> , \RAM<48><2> , \RAM<48><1> , \RAM<48><0> , \RAM<47><31> ,
         \RAM<47><30> , \RAM<47><29> , \RAM<47><28> , \RAM<47><27> ,
         \RAM<47><26> , \RAM<47><25> , \RAM<47><24> , \RAM<47><23> ,
         \RAM<47><22> , \RAM<47><21> , \RAM<47><20> , \RAM<47><19> ,
         \RAM<47><18> , \RAM<47><17> , \RAM<47><16> , \RAM<47><15> ,
         \RAM<47><14> , \RAM<47><13> , \RAM<47><12> , \RAM<47><11> ,
         \RAM<47><10> , \RAM<47><9> , \RAM<47><8> , \RAM<47><7> , \RAM<47><6> ,
         \RAM<47><5> , \RAM<47><4> , \RAM<47><3> , \RAM<47><2> , \RAM<47><1> ,
         \RAM<47><0> , \RAM<46><31> , \RAM<46><30> , \RAM<46><29> ,
         \RAM<46><28> , \RAM<46><27> , \RAM<46><26> , \RAM<46><25> ,
         \RAM<46><24> , \RAM<46><23> , \RAM<46><22> , \RAM<46><21> ,
         \RAM<46><20> , \RAM<46><19> , \RAM<46><18> , \RAM<46><17> ,
         \RAM<46><16> , \RAM<46><15> , \RAM<46><14> , \RAM<46><13> ,
         \RAM<46><12> , \RAM<46><11> , \RAM<46><10> , \RAM<46><9> ,
         \RAM<46><8> , \RAM<46><7> , \RAM<46><6> , \RAM<46><5> , \RAM<46><4> ,
         \RAM<46><3> , \RAM<46><2> , \RAM<46><1> , \RAM<46><0> , \RAM<45><31> ,
         \RAM<45><30> , \RAM<45><29> , \RAM<45><28> , \RAM<45><27> ,
         \RAM<45><26> , \RAM<45><25> , \RAM<45><24> , \RAM<45><23> ,
         \RAM<45><22> , \RAM<45><21> , \RAM<45><20> , \RAM<45><19> ,
         \RAM<45><18> , \RAM<45><17> , \RAM<45><16> , \RAM<45><15> ,
         \RAM<45><14> , \RAM<45><13> , \RAM<45><12> , \RAM<45><11> ,
         \RAM<45><10> , \RAM<45><9> , \RAM<45><8> , \RAM<45><7> , \RAM<45><6> ,
         \RAM<45><5> , \RAM<45><4> , \RAM<45><3> , \RAM<45><2> , \RAM<45><1> ,
         \RAM<45><0> , \RAM<44><31> , \RAM<44><30> , \RAM<44><29> ,
         \RAM<44><28> , \RAM<44><27> , \RAM<44><26> , \RAM<44><25> ,
         \RAM<44><24> , \RAM<44><23> , \RAM<44><22> , \RAM<44><21> ,
         \RAM<44><20> , \RAM<44><19> , \RAM<44><18> , \RAM<44><17> ,
         \RAM<44><16> , \RAM<44><15> , \RAM<44><14> , \RAM<44><13> ,
         \RAM<44><12> , \RAM<44><11> , \RAM<44><10> , \RAM<44><9> ,
         \RAM<44><8> , \RAM<44><7> , \RAM<44><6> , \RAM<44><5> , \RAM<44><4> ,
         \RAM<44><3> , \RAM<44><2> , \RAM<44><1> , \RAM<44><0> , \RAM<43><31> ,
         \RAM<43><30> , \RAM<43><29> , \RAM<43><28> , \RAM<43><27> ,
         \RAM<43><26> , \RAM<43><25> , \RAM<43><24> , \RAM<43><23> ,
         \RAM<43><22> , \RAM<43><21> , \RAM<43><20> , \RAM<43><19> ,
         \RAM<43><18> , \RAM<43><17> , \RAM<43><16> , \RAM<43><15> ,
         \RAM<43><14> , \RAM<43><13> , \RAM<43><12> , \RAM<43><11> ,
         \RAM<43><10> , \RAM<43><9> , \RAM<43><8> , \RAM<43><7> , \RAM<43><6> ,
         \RAM<43><5> , \RAM<43><4> , \RAM<43><3> , \RAM<43><2> , \RAM<43><1> ,
         \RAM<43><0> , \RAM<42><31> , \RAM<42><30> , \RAM<42><29> ,
         \RAM<42><28> , \RAM<42><27> , \RAM<42><26> , \RAM<42><25> ,
         \RAM<42><24> , \RAM<42><23> , \RAM<42><22> , \RAM<42><21> ,
         \RAM<42><20> , \RAM<42><19> , \RAM<42><18> , \RAM<42><17> ,
         \RAM<42><16> , \RAM<42><15> , \RAM<42><14> , \RAM<42><13> ,
         \RAM<42><12> , \RAM<42><11> , \RAM<42><10> , \RAM<42><9> ,
         \RAM<42><8> , \RAM<42><7> , \RAM<42><6> , \RAM<42><5> , \RAM<42><4> ,
         \RAM<42><3> , \RAM<42><2> , \RAM<42><1> , \RAM<42><0> , \RAM<41><31> ,
         \RAM<41><30> , \RAM<41><29> , \RAM<41><28> , \RAM<41><27> ,
         \RAM<41><26> , \RAM<41><25> , \RAM<41><24> , \RAM<41><23> ,
         \RAM<41><22> , \RAM<41><21> , \RAM<41><20> , \RAM<41><19> ,
         \RAM<41><18> , \RAM<41><17> , \RAM<41><16> , \RAM<41><15> ,
         \RAM<41><14> , \RAM<41><13> , \RAM<41><12> , \RAM<41><11> ,
         \RAM<41><10> , \RAM<41><9> , \RAM<41><8> , \RAM<41><7> , \RAM<41><6> ,
         \RAM<41><5> , \RAM<41><4> , \RAM<41><3> , \RAM<41><2> , \RAM<41><1> ,
         \RAM<41><0> , \RAM<40><31> , \RAM<40><30> , \RAM<40><29> ,
         \RAM<40><28> , \RAM<40><27> , \RAM<40><26> , \RAM<40><25> ,
         \RAM<40><24> , \RAM<40><23> , \RAM<40><22> , \RAM<40><21> ,
         \RAM<40><20> , \RAM<40><19> , \RAM<40><18> , \RAM<40><17> ,
         \RAM<40><16> , \RAM<40><15> , \RAM<40><14> , \RAM<40><13> ,
         \RAM<40><12> , \RAM<40><11> , \RAM<40><10> , \RAM<40><9> ,
         \RAM<40><8> , \RAM<40><7> , \RAM<40><6> , \RAM<40><5> , \RAM<40><4> ,
         \RAM<40><3> , \RAM<40><2> , \RAM<40><1> , \RAM<40><0> , \RAM<39><31> ,
         \RAM<39><30> , \RAM<39><29> , \RAM<39><28> , \RAM<39><27> ,
         \RAM<39><26> , \RAM<39><25> , \RAM<39><24> , \RAM<39><23> ,
         \RAM<39><22> , \RAM<39><21> , \RAM<39><20> , \RAM<39><19> ,
         \RAM<39><18> , \RAM<39><17> , \RAM<39><16> , \RAM<39><15> ,
         \RAM<39><14> , \RAM<39><13> , \RAM<39><12> , \RAM<39><11> ,
         \RAM<39><10> , \RAM<39><9> , \RAM<39><8> , \RAM<39><7> , \RAM<39><6> ,
         \RAM<39><5> , \RAM<39><4> , \RAM<39><3> , \RAM<39><2> , \RAM<39><1> ,
         \RAM<39><0> , \RAM<38><31> , \RAM<38><30> , \RAM<38><29> ,
         \RAM<38><28> , \RAM<38><27> , \RAM<38><26> , \RAM<38><25> ,
         \RAM<38><24> , \RAM<38><23> , \RAM<38><22> , \RAM<38><21> ,
         \RAM<38><20> , \RAM<38><19> , \RAM<38><18> , \RAM<38><17> ,
         \RAM<38><16> , \RAM<38><15> , \RAM<38><14> , \RAM<38><13> ,
         \RAM<38><12> , \RAM<38><11> , \RAM<38><10> , \RAM<38><9> ,
         \RAM<38><8> , \RAM<38><7> , \RAM<38><6> , \RAM<38><5> , \RAM<38><4> ,
         \RAM<38><3> , \RAM<38><2> , \RAM<38><1> , \RAM<38><0> , \RAM<37><31> ,
         \RAM<37><30> , \RAM<37><29> , \RAM<37><28> , \RAM<37><27> ,
         \RAM<37><26> , \RAM<37><25> , \RAM<37><24> , \RAM<37><23> ,
         \RAM<37><22> , \RAM<37><21> , \RAM<37><20> , \RAM<37><19> ,
         \RAM<37><18> , \RAM<37><17> , \RAM<37><16> , \RAM<37><15> ,
         \RAM<37><14> , \RAM<37><13> , \RAM<37><12> , \RAM<37><11> ,
         \RAM<37><10> , \RAM<37><9> , \RAM<37><8> , \RAM<37><7> , \RAM<37><6> ,
         \RAM<37><5> , \RAM<37><4> , \RAM<37><3> , \RAM<37><2> , \RAM<37><1> ,
         \RAM<37><0> , \RAM<36><31> , \RAM<36><30> , \RAM<36><29> ,
         \RAM<36><28> , \RAM<36><27> , \RAM<36><26> , \RAM<36><25> ,
         \RAM<36><24> , \RAM<36><23> , \RAM<36><22> , \RAM<36><21> ,
         \RAM<36><20> , \RAM<36><19> , \RAM<36><18> , \RAM<36><17> ,
         \RAM<36><16> , \RAM<36><15> , \RAM<36><14> , \RAM<36><13> ,
         \RAM<36><12> , \RAM<36><11> , \RAM<36><10> , \RAM<36><9> ,
         \RAM<36><8> , \RAM<36><7> , \RAM<36><6> , \RAM<36><5> , \RAM<36><4> ,
         \RAM<36><3> , \RAM<36><2> , \RAM<36><1> , \RAM<36><0> , \RAM<35><31> ,
         \RAM<35><30> , \RAM<35><29> , \RAM<35><28> , \RAM<35><27> ,
         \RAM<35><26> , \RAM<35><25> , \RAM<35><24> , \RAM<35><23> ,
         \RAM<35><22> , \RAM<35><21> , \RAM<35><20> , \RAM<35><19> ,
         \RAM<35><18> , \RAM<35><17> , \RAM<35><16> , \RAM<35><15> ,
         \RAM<35><14> , \RAM<35><13> , \RAM<35><12> , \RAM<35><11> ,
         \RAM<35><10> , \RAM<35><9> , \RAM<35><8> , \RAM<35><7> , \RAM<35><6> ,
         \RAM<35><5> , \RAM<35><4> , \RAM<35><3> , \RAM<35><2> , \RAM<35><1> ,
         \RAM<35><0> , \RAM<34><31> , \RAM<34><30> , \RAM<34><29> ,
         \RAM<34><28> , \RAM<34><27> , \RAM<34><26> , \RAM<34><25> ,
         \RAM<34><24> , \RAM<34><23> , \RAM<34><22> , \RAM<34><21> ,
         \RAM<34><20> , \RAM<34><19> , \RAM<34><18> , \RAM<34><17> ,
         \RAM<34><16> , \RAM<34><15> , \RAM<34><14> , \RAM<34><13> ,
         \RAM<34><12> , \RAM<34><11> , \RAM<34><10> , \RAM<34><9> ,
         \RAM<34><8> , \RAM<34><7> , \RAM<34><6> , \RAM<34><5> , \RAM<34><4> ,
         \RAM<34><3> , \RAM<34><2> , \RAM<34><1> , \RAM<34><0> , \RAM<33><31> ,
         \RAM<33><30> , \RAM<33><29> , \RAM<33><28> , \RAM<33><27> ,
         \RAM<33><26> , \RAM<33><25> , \RAM<33><24> , \RAM<33><23> ,
         \RAM<33><22> , \RAM<33><21> , \RAM<33><20> , \RAM<33><19> ,
         \RAM<33><18> , \RAM<33><17> , \RAM<33><16> , \RAM<33><15> ,
         \RAM<33><14> , \RAM<33><13> , \RAM<33><12> , \RAM<33><11> ,
         \RAM<33><10> , \RAM<33><9> , \RAM<33><8> , \RAM<33><7> , \RAM<33><6> ,
         \RAM<33><5> , \RAM<33><4> , \RAM<33><3> , \RAM<33><2> , \RAM<33><1> ,
         \RAM<33><0> , \RAM<32><31> , \RAM<32><30> , \RAM<32><29> ,
         \RAM<32><28> , \RAM<32><27> , \RAM<32><26> , \RAM<32><25> ,
         \RAM<32><24> , \RAM<32><23> , \RAM<32><22> , \RAM<32><21> ,
         \RAM<32><20> , \RAM<32><19> , \RAM<32><18> , \RAM<32><17> ,
         \RAM<32><16> , \RAM<32><15> , \RAM<32><14> , \RAM<32><13> ,
         \RAM<32><12> , \RAM<32><11> , \RAM<32><10> , \RAM<32><9> ,
         \RAM<32><8> , \RAM<32><7> , \RAM<32><6> , \RAM<32><5> , \RAM<32><4> ,
         \RAM<32><3> , \RAM<32><2> , \RAM<32><1> , \RAM<32><0> , \RAM<31><31> ,
         \RAM<31><30> , \RAM<31><29> , \RAM<31><28> , \RAM<31><27> ,
         \RAM<31><26> , \RAM<31><25> , \RAM<31><24> , \RAM<31><23> ,
         \RAM<31><22> , \RAM<31><21> , \RAM<31><20> , \RAM<31><19> ,
         \RAM<31><18> , \RAM<31><17> , \RAM<31><16> , \RAM<31><15> ,
         \RAM<31><14> , \RAM<31><13> , \RAM<31><12> , \RAM<31><11> ,
         \RAM<31><10> , \RAM<31><9> , \RAM<31><8> , \RAM<31><7> , \RAM<31><6> ,
         \RAM<31><5> , \RAM<31><4> , \RAM<31><3> , \RAM<31><2> , \RAM<31><1> ,
         \RAM<31><0> , \RAM<30><31> , \RAM<30><30> , \RAM<30><29> ,
         \RAM<30><28> , \RAM<30><27> , \RAM<30><26> , \RAM<30><25> ,
         \RAM<30><24> , \RAM<30><23> , \RAM<30><22> , \RAM<30><21> ,
         \RAM<30><20> , \RAM<30><19> , \RAM<30><18> , \RAM<30><17> ,
         \RAM<30><16> , \RAM<30><15> , \RAM<30><14> , \RAM<30><13> ,
         \RAM<30><12> , \RAM<30><11> , \RAM<30><10> , \RAM<30><9> ,
         \RAM<30><8> , \RAM<30><7> , \RAM<30><6> , \RAM<30><5> , \RAM<30><4> ,
         \RAM<30><3> , \RAM<30><2> , \RAM<30><1> , \RAM<30><0> , \RAM<29><31> ,
         \RAM<29><30> , \RAM<29><29> , \RAM<29><28> , \RAM<29><27> ,
         \RAM<29><26> , \RAM<29><25> , \RAM<29><24> , \RAM<29><23> ,
         \RAM<29><22> , \RAM<29><21> , \RAM<29><20> , \RAM<29><19> ,
         \RAM<29><18> , \RAM<29><17> , \RAM<29><16> , \RAM<29><15> ,
         \RAM<29><14> , \RAM<29><13> , \RAM<29><12> , \RAM<29><11> ,
         \RAM<29><10> , \RAM<29><9> , \RAM<29><8> , \RAM<29><7> , \RAM<29><6> ,
         \RAM<29><5> , \RAM<29><4> , \RAM<29><3> , \RAM<29><2> , \RAM<29><1> ,
         \RAM<29><0> , \RAM<28><31> , \RAM<28><30> , \RAM<28><29> ,
         \RAM<28><28> , \RAM<28><27> , \RAM<28><26> , \RAM<28><25> ,
         \RAM<28><24> , \RAM<28><23> , \RAM<28><22> , \RAM<28><21> ,
         \RAM<28><20> , \RAM<28><19> , \RAM<28><18> , \RAM<28><17> ,
         \RAM<28><16> , \RAM<28><15> , \RAM<28><14> , \RAM<28><13> ,
         \RAM<28><12> , \RAM<28><11> , \RAM<28><10> , \RAM<28><9> ,
         \RAM<28><8> , \RAM<28><7> , \RAM<28><6> , \RAM<28><5> , \RAM<28><4> ,
         \RAM<28><3> , \RAM<28><2> , \RAM<28><1> , \RAM<28><0> , \RAM<27><31> ,
         \RAM<27><30> , \RAM<27><29> , \RAM<27><28> , \RAM<27><27> ,
         \RAM<27><26> , \RAM<27><25> , \RAM<27><24> , \RAM<27><23> ,
         \RAM<27><22> , \RAM<27><21> , \RAM<27><20> , \RAM<27><19> ,
         \RAM<27><18> , \RAM<27><17> , \RAM<27><16> , \RAM<27><15> ,
         \RAM<27><14> , \RAM<27><13> , \RAM<27><12> , \RAM<27><11> ,
         \RAM<27><10> , \RAM<27><9> , \RAM<27><8> , \RAM<27><7> , \RAM<27><6> ,
         \RAM<27><5> , \RAM<27><4> , \RAM<27><3> , \RAM<27><2> , \RAM<27><1> ,
         \RAM<27><0> , \RAM<26><31> , \RAM<26><30> , \RAM<26><29> ,
         \RAM<26><28> , \RAM<26><27> , \RAM<26><26> , \RAM<26><25> ,
         \RAM<26><24> , \RAM<26><23> , \RAM<26><22> , \RAM<26><21> ,
         \RAM<26><20> , \RAM<26><19> , \RAM<26><18> , \RAM<26><17> ,
         \RAM<26><16> , \RAM<26><15> , \RAM<26><14> , \RAM<26><13> ,
         \RAM<26><12> , \RAM<26><11> , \RAM<26><10> , \RAM<26><9> ,
         \RAM<26><8> , \RAM<26><7> , \RAM<26><6> , \RAM<26><5> , \RAM<26><4> ,
         \RAM<26><3> , \RAM<26><2> , \RAM<26><1> , \RAM<26><0> , \RAM<25><31> ,
         \RAM<25><30> , \RAM<25><29> , \RAM<25><28> , \RAM<25><27> ,
         \RAM<25><26> , \RAM<25><25> , \RAM<25><24> , \RAM<25><23> ,
         \RAM<25><22> , \RAM<25><21> , \RAM<25><20> , \RAM<25><19> ,
         \RAM<25><18> , \RAM<25><17> , \RAM<25><16> , \RAM<25><15> ,
         \RAM<25><14> , \RAM<25><13> , \RAM<25><12> , \RAM<25><11> ,
         \RAM<25><10> , \RAM<25><9> , \RAM<25><8> , \RAM<25><7> , \RAM<25><6> ,
         \RAM<25><5> , \RAM<25><4> , \RAM<25><3> , \RAM<25><2> , \RAM<25><1> ,
         \RAM<25><0> , \RAM<24><31> , \RAM<24><30> , \RAM<24><29> ,
         \RAM<24><28> , \RAM<24><27> , \RAM<24><26> , \RAM<24><25> ,
         \RAM<24><24> , \RAM<24><23> , \RAM<24><22> , \RAM<24><21> ,
         \RAM<24><20> , \RAM<24><19> , \RAM<24><18> , \RAM<24><17> ,
         \RAM<24><16> , \RAM<24><15> , \RAM<24><14> , \RAM<24><13> ,
         \RAM<24><12> , \RAM<24><11> , \RAM<24><10> , \RAM<24><9> ,
         \RAM<24><8> , \RAM<24><7> , \RAM<24><6> , \RAM<24><5> , \RAM<24><4> ,
         \RAM<24><3> , \RAM<24><2> , \RAM<24><1> , \RAM<24><0> , \RAM<23><31> ,
         \RAM<23><30> , \RAM<23><29> , \RAM<23><28> , \RAM<23><27> ,
         \RAM<23><26> , \RAM<23><25> , \RAM<23><24> , \RAM<23><23> ,
         \RAM<23><22> , \RAM<23><21> , \RAM<23><20> , \RAM<23><19> ,
         \RAM<23><18> , \RAM<23><17> , \RAM<23><16> , \RAM<23><15> ,
         \RAM<23><14> , \RAM<23><13> , \RAM<23><12> , \RAM<23><11> ,
         \RAM<23><10> , \RAM<23><9> , \RAM<23><8> , \RAM<23><7> , \RAM<23><6> ,
         \RAM<23><5> , \RAM<23><4> , \RAM<23><3> , \RAM<23><2> , \RAM<23><1> ,
         \RAM<23><0> , \RAM<22><31> , \RAM<22><30> , \RAM<22><29> ,
         \RAM<22><28> , \RAM<22><27> , \RAM<22><26> , \RAM<22><25> ,
         \RAM<22><24> , \RAM<22><23> , \RAM<22><22> , \RAM<22><21> ,
         \RAM<22><20> , \RAM<22><19> , \RAM<22><18> , \RAM<22><17> ,
         \RAM<22><16> , \RAM<22><15> , \RAM<22><14> , \RAM<22><13> ,
         \RAM<22><12> , \RAM<22><11> , \RAM<22><10> , \RAM<22><9> ,
         \RAM<22><8> , \RAM<22><7> , \RAM<22><6> , \RAM<22><5> , \RAM<22><4> ,
         \RAM<22><3> , \RAM<22><2> , \RAM<22><1> , \RAM<22><0> , \RAM<21><31> ,
         \RAM<21><30> , \RAM<21><29> , \RAM<21><28> , \RAM<21><27> ,
         \RAM<21><26> , \RAM<21><25> , \RAM<21><24> , \RAM<21><23> ,
         \RAM<21><22> , \RAM<21><21> , \RAM<21><20> , \RAM<21><19> ,
         \RAM<21><18> , \RAM<21><17> , \RAM<21><16> , \RAM<21><15> ,
         \RAM<21><14> , \RAM<21><13> , \RAM<21><12> , \RAM<21><11> ,
         \RAM<21><10> , \RAM<21><9> , \RAM<21><8> , \RAM<21><7> , \RAM<21><6> ,
         \RAM<21><5> , \RAM<21><4> , \RAM<21><3> , \RAM<21><2> , \RAM<21><1> ,
         \RAM<21><0> , \RAM<20><31> , \RAM<20><30> , \RAM<20><29> ,
         \RAM<20><28> , \RAM<20><27> , \RAM<20><26> , \RAM<20><25> ,
         \RAM<20><24> , \RAM<20><23> , \RAM<20><22> , \RAM<20><21> ,
         \RAM<20><20> , \RAM<20><19> , \RAM<20><18> , \RAM<20><17> ,
         \RAM<20><16> , \RAM<20><15> , \RAM<20><14> , \RAM<20><13> ,
         \RAM<20><12> , \RAM<20><11> , \RAM<20><10> , \RAM<20><9> ,
         \RAM<20><8> , \RAM<20><7> , \RAM<20><6> , \RAM<20><5> , \RAM<20><4> ,
         \RAM<20><3> , \RAM<20><2> , \RAM<20><1> , \RAM<20><0> , \RAM<19><31> ,
         \RAM<19><30> , \RAM<19><29> , \RAM<19><28> , \RAM<19><27> ,
         \RAM<19><26> , \RAM<19><25> , \RAM<19><24> , \RAM<19><23> ,
         \RAM<19><22> , \RAM<19><21> , \RAM<19><20> , \RAM<19><19> ,
         \RAM<19><18> , \RAM<19><17> , \RAM<19><16> , \RAM<19><15> ,
         \RAM<19><14> , \RAM<19><13> , \RAM<19><12> , \RAM<19><11> ,
         \RAM<19><10> , \RAM<19><9> , \RAM<19><8> , \RAM<19><7> , \RAM<19><6> ,
         \RAM<19><5> , \RAM<19><4> , \RAM<19><3> , \RAM<19><2> , \RAM<19><1> ,
         \RAM<19><0> , \RAM<18><31> , \RAM<18><30> , \RAM<18><29> ,
         \RAM<18><28> , \RAM<18><27> , \RAM<18><26> , \RAM<18><25> ,
         \RAM<18><24> , \RAM<18><23> , \RAM<18><22> , \RAM<18><21> ,
         \RAM<18><20> , \RAM<18><19> , \RAM<18><18> , \RAM<18><17> ,
         \RAM<18><16> , \RAM<18><15> , \RAM<18><14> , \RAM<18><13> ,
         \RAM<18><12> , \RAM<18><11> , \RAM<18><10> , \RAM<18><9> ,
         \RAM<18><8> , \RAM<18><7> , \RAM<18><6> , \RAM<18><5> , \RAM<18><4> ,
         \RAM<18><3> , \RAM<18><2> , \RAM<18><1> , \RAM<18><0> , \RAM<17><31> ,
         \RAM<17><30> , \RAM<17><29> , \RAM<17><28> , \RAM<17><27> ,
         \RAM<17><26> , \RAM<17><25> , \RAM<17><24> , \RAM<17><23> ,
         \RAM<17><22> , \RAM<17><21> , \RAM<17><20> , \RAM<17><19> ,
         \RAM<17><18> , \RAM<17><17> , \RAM<17><16> , \RAM<17><15> ,
         \RAM<17><14> , \RAM<17><13> , \RAM<17><12> , \RAM<17><11> ,
         \RAM<17><10> , \RAM<17><9> , \RAM<17><8> , \RAM<17><7> , \RAM<17><6> ,
         \RAM<17><5> , \RAM<17><4> , \RAM<17><3> , \RAM<17><2> , \RAM<17><1> ,
         \RAM<17><0> , \RAM<16><31> , \RAM<16><30> , \RAM<16><29> ,
         \RAM<16><28> , \RAM<16><27> , \RAM<16><26> , \RAM<16><25> ,
         \RAM<16><24> , \RAM<16><23> , \RAM<16><22> , \RAM<16><21> ,
         \RAM<16><20> , \RAM<16><19> , \RAM<16><18> , \RAM<16><17> ,
         \RAM<16><16> , \RAM<16><15> , \RAM<16><14> , \RAM<16><13> ,
         \RAM<16><12> , \RAM<16><11> , \RAM<16><10> , \RAM<16><9> ,
         \RAM<16><8> , \RAM<16><7> , \RAM<16><6> , \RAM<16><5> , \RAM<16><4> ,
         \RAM<16><3> , \RAM<16><2> , \RAM<16><1> , \RAM<16><0> , \RAM<15><31> ,
         \RAM<15><30> , \RAM<15><29> , \RAM<15><28> , \RAM<15><27> ,
         \RAM<15><26> , \RAM<15><25> , \RAM<15><24> , \RAM<15><23> ,
         \RAM<15><22> , \RAM<15><21> , \RAM<15><20> , \RAM<15><19> ,
         \RAM<15><18> , \RAM<15><17> , \RAM<15><16> , \RAM<15><15> ,
         \RAM<15><14> , \RAM<15><13> , \RAM<15><12> , \RAM<15><11> ,
         \RAM<15><10> , \RAM<15><9> , \RAM<15><8> , \RAM<15><7> , \RAM<15><6> ,
         \RAM<15><5> , \RAM<15><4> , \RAM<15><3> , \RAM<15><2> , \RAM<15><1> ,
         \RAM<15><0> , \RAM<14><31> , \RAM<14><30> , \RAM<14><29> ,
         \RAM<14><28> , \RAM<14><27> , \RAM<14><26> , \RAM<14><25> ,
         \RAM<14><24> , \RAM<14><23> , \RAM<14><22> , \RAM<14><21> ,
         \RAM<14><20> , \RAM<14><19> , \RAM<14><18> , \RAM<14><17> ,
         \RAM<14><16> , \RAM<14><15> , \RAM<14><14> , \RAM<14><13> ,
         \RAM<14><12> , \RAM<14><11> , \RAM<14><10> , \RAM<14><9> ,
         \RAM<14><8> , \RAM<14><7> , \RAM<14><6> , \RAM<14><5> , \RAM<14><4> ,
         \RAM<14><3> , \RAM<14><2> , \RAM<14><1> , \RAM<14><0> , \RAM<13><31> ,
         \RAM<13><30> , \RAM<13><29> , \RAM<13><28> , \RAM<13><27> ,
         \RAM<13><26> , \RAM<13><25> , \RAM<13><24> , \RAM<13><23> ,
         \RAM<13><22> , \RAM<13><21> , \RAM<13><20> , \RAM<13><19> ,
         \RAM<13><18> , \RAM<13><17> , \RAM<13><16> , \RAM<13><15> ,
         \RAM<13><14> , \RAM<13><13> , \RAM<13><12> , \RAM<13><11> ,
         \RAM<13><10> , \RAM<13><9> , \RAM<13><8> , \RAM<13><7> , \RAM<13><6> ,
         \RAM<13><5> , \RAM<13><4> , \RAM<13><3> , \RAM<13><2> , \RAM<13><1> ,
         \RAM<13><0> , \RAM<12><31> , \RAM<12><30> , \RAM<12><29> ,
         \RAM<12><28> , \RAM<12><27> , \RAM<12><26> , \RAM<12><25> ,
         \RAM<12><24> , \RAM<12><23> , \RAM<12><22> , \RAM<12><21> ,
         \RAM<12><20> , \RAM<12><19> , \RAM<12><18> , \RAM<12><17> ,
         \RAM<12><16> , \RAM<12><15> , \RAM<12><14> , \RAM<12><13> ,
         \RAM<12><12> , \RAM<12><11> , \RAM<12><10> , \RAM<12><9> ,
         \RAM<12><8> , \RAM<12><7> , \RAM<12><6> , \RAM<12><5> , \RAM<12><4> ,
         \RAM<12><3> , \RAM<12><2> , \RAM<12><1> , \RAM<12><0> , \RAM<11><31> ,
         \RAM<11><30> , \RAM<11><29> , \RAM<11><28> , \RAM<11><27> ,
         \RAM<11><26> , \RAM<11><25> , \RAM<11><24> , \RAM<11><23> ,
         \RAM<11><22> , \RAM<11><21> , \RAM<11><20> , \RAM<11><19> ,
         \RAM<11><18> , \RAM<11><17> , \RAM<11><16> , \RAM<11><15> ,
         \RAM<11><14> , \RAM<11><13> , \RAM<11><12> , \RAM<11><11> ,
         \RAM<11><10> , \RAM<11><9> , \RAM<11><8> , \RAM<11><7> , \RAM<11><6> ,
         \RAM<11><5> , \RAM<11><4> , \RAM<11><3> , \RAM<11><2> , \RAM<11><1> ,
         \RAM<11><0> , \RAM<10><31> , \RAM<10><30> , \RAM<10><29> ,
         \RAM<10><28> , \RAM<10><27> , \RAM<10><26> , \RAM<10><25> ,
         \RAM<10><24> , \RAM<10><23> , \RAM<10><22> , \RAM<10><21> ,
         \RAM<10><20> , \RAM<10><19> , \RAM<10><18> , \RAM<10><17> ,
         \RAM<10><16> , \RAM<10><15> , \RAM<10><14> , \RAM<10><13> ,
         \RAM<10><12> , \RAM<10><11> , \RAM<10><10> , \RAM<10><9> ,
         \RAM<10><8> , \RAM<10><7> , \RAM<10><6> , \RAM<10><5> , \RAM<10><4> ,
         \RAM<10><3> , \RAM<10><2> , \RAM<10><1> , \RAM<10><0> , \RAM<9><31> ,
         \RAM<9><30> , \RAM<9><29> , \RAM<9><28> , \RAM<9><27> , \RAM<9><26> ,
         \RAM<9><25> , \RAM<9><24> , \RAM<9><23> , \RAM<9><22> , \RAM<9><21> ,
         \RAM<9><20> , \RAM<9><19> , \RAM<9><18> , \RAM<9><17> , \RAM<9><16> ,
         \RAM<9><15> , \RAM<9><14> , \RAM<9><13> , \RAM<9><12> , \RAM<9><11> ,
         \RAM<9><10> , \RAM<9><9> , \RAM<9><8> , \RAM<9><7> , \RAM<9><6> ,
         \RAM<9><5> , \RAM<9><4> , \RAM<9><3> , \RAM<9><2> , \RAM<9><1> ,
         \RAM<9><0> , \RAM<8><31> , \RAM<8><30> , \RAM<8><29> , \RAM<8><28> ,
         \RAM<8><27> , \RAM<8><26> , \RAM<8><25> , \RAM<8><24> , \RAM<8><23> ,
         \RAM<8><22> , \RAM<8><21> , \RAM<8><20> , \RAM<8><19> , \RAM<8><18> ,
         \RAM<8><17> , \RAM<8><16> , \RAM<8><15> , \RAM<8><14> , \RAM<8><13> ,
         \RAM<8><12> , \RAM<8><11> , \RAM<8><10> , \RAM<8><9> , \RAM<8><8> ,
         \RAM<8><7> , \RAM<8><6> , \RAM<8><5> , \RAM<8><4> , \RAM<8><3> ,
         \RAM<8><2> , \RAM<8><1> , \RAM<8><0> , \RAM<7><31> , \RAM<7><30> ,
         \RAM<7><29> , \RAM<7><28> , \RAM<7><27> , \RAM<7><26> , \RAM<7><25> ,
         \RAM<7><24> , \RAM<7><23> , \RAM<7><22> , \RAM<7><21> , \RAM<7><20> ,
         \RAM<7><19> , \RAM<7><18> , \RAM<7><17> , \RAM<7><16> , \RAM<7><15> ,
         \RAM<7><14> , \RAM<7><13> , \RAM<7><12> , \RAM<7><11> , \RAM<7><10> ,
         \RAM<7><9> , \RAM<7><8> , \RAM<7><7> , \RAM<7><6> , \RAM<7><5> ,
         \RAM<7><4> , \RAM<7><3> , \RAM<7><2> , \RAM<7><1> , \RAM<7><0> ,
         \RAM<6><31> , \RAM<6><30> , \RAM<6><29> , \RAM<6><28> , \RAM<6><27> ,
         \RAM<6><26> , \RAM<6><25> , \RAM<6><24> , \RAM<6><23> , \RAM<6><22> ,
         \RAM<6><21> , \RAM<6><20> , \RAM<6><19> , \RAM<6><18> , \RAM<6><17> ,
         \RAM<6><16> , \RAM<6><15> , \RAM<6><14> , \RAM<6><13> , \RAM<6><12> ,
         \RAM<6><11> , \RAM<6><10> , \RAM<6><9> , \RAM<6><8> , \RAM<6><7> ,
         \RAM<6><6> , \RAM<6><5> , \RAM<6><4> , \RAM<6><3> , \RAM<6><2> ,
         \RAM<6><1> , \RAM<6><0> , \RAM<5><31> , \RAM<5><30> , \RAM<5><29> ,
         \RAM<5><28> , \RAM<5><27> , \RAM<5><26> , \RAM<5><25> , \RAM<5><24> ,
         \RAM<5><23> , \RAM<5><22> , \RAM<5><21> , \RAM<5><20> , \RAM<5><19> ,
         \RAM<5><18> , \RAM<5><17> , \RAM<5><16> , \RAM<5><15> , \RAM<5><14> ,
         \RAM<5><13> , \RAM<5><12> , \RAM<5><11> , \RAM<5><10> , \RAM<5><9> ,
         \RAM<5><8> , \RAM<5><7> , \RAM<5><6> , \RAM<5><5> , \RAM<5><4> ,
         \RAM<5><3> , \RAM<5><2> , \RAM<5><1> , \RAM<5><0> , \RAM<4><31> ,
         \RAM<4><30> , \RAM<4><29> , \RAM<4><28> , \RAM<4><27> , \RAM<4><26> ,
         \RAM<4><25> , \RAM<4><24> , \RAM<4><23> , \RAM<4><22> , \RAM<4><21> ,
         \RAM<4><20> , \RAM<4><19> , \RAM<4><18> , \RAM<4><17> , \RAM<4><16> ,
         \RAM<4><15> , \RAM<4><14> , \RAM<4><13> , \RAM<4><12> , \RAM<4><11> ,
         \RAM<4><10> , \RAM<4><9> , \RAM<4><8> , \RAM<4><7> , \RAM<4><6> ,
         \RAM<4><5> , \RAM<4><4> , \RAM<4><3> , \RAM<4><2> , \RAM<4><1> ,
         \RAM<4><0> , \RAM<3><31> , \RAM<3><30> , \RAM<3><29> , \RAM<3><28> ,
         \RAM<3><27> , \RAM<3><26> , \RAM<3><25> , \RAM<3><24> , \RAM<3><23> ,
         \RAM<3><22> , \RAM<3><21> , \RAM<3><20> , \RAM<3><19> , \RAM<3><18> ,
         \RAM<3><17> , \RAM<3><16> , \RAM<3><15> , \RAM<3><14> , \RAM<3><13> ,
         \RAM<3><12> , \RAM<3><11> , \RAM<3><10> , \RAM<3><9> , \RAM<3><8> ,
         \RAM<3><7> , \RAM<3><6> , \RAM<3><5> , \RAM<3><4> , \RAM<3><3> ,
         \RAM<3><2> , \RAM<3><1> , \RAM<3><0> , \RAM<2><31> , \RAM<2><30> ,
         \RAM<2><29> , \RAM<2><28> , \RAM<2><27> , \RAM<2><26> , \RAM<2><25> ,
         \RAM<2><24> , \RAM<2><23> , \RAM<2><22> , \RAM<2><21> , \RAM<2><20> ,
         \RAM<2><19> , \RAM<2><18> , \RAM<2><17> , \RAM<2><16> , \RAM<2><15> ,
         \RAM<2><14> , \RAM<2><13> , \RAM<2><12> , \RAM<2><11> , \RAM<2><10> ,
         \RAM<2><9> , \RAM<2><8> , \RAM<2><7> , \RAM<2><6> , \RAM<2><5> ,
         \RAM<2><4> , \RAM<2><3> , \RAM<2><2> , \RAM<2><1> , \RAM<2><0> ,
         \RAM<1><31> , \RAM<1><30> , \RAM<1><29> , \RAM<1><28> , \RAM<1><27> ,
         \RAM<1><26> , \RAM<1><25> , \RAM<1><24> , \RAM<1><23> , \RAM<1><22> ,
         \RAM<1><21> , \RAM<1><20> , \RAM<1><19> , \RAM<1><18> , \RAM<1><17> ,
         \RAM<1><16> , \RAM<1><15> , \RAM<1><14> , \RAM<1><13> , \RAM<1><12> ,
         \RAM<1><11> , \RAM<1><10> , \RAM<1><9> , \RAM<1><8> , \RAM<1><7> ,
         \RAM<1><6> , \RAM<1><5> , \RAM<1><4> , \RAM<1><3> , \RAM<1><2> ,
         \RAM<1><1> , \RAM<1><0> , \RAM<0><31> , \RAM<0><30> , \RAM<0><29> ,
         \RAM<0><28> , \RAM<0><27> , \RAM<0><26> , \RAM<0><25> , \RAM<0><24> ,
         \RAM<0><23> , \RAM<0><22> , \RAM<0><21> , \RAM<0><20> , \RAM<0><19> ,
         \RAM<0><18> , \RAM<0><17> , \RAM<0><16> , \RAM<0><15> , \RAM<0><14> ,
         \RAM<0><13> , \RAM<0><12> , \RAM<0><11> , \RAM<0><10> , \RAM<0><9> ,
         \RAM<0><8> , \RAM<0><7> , \RAM<0><6> , \RAM<0><5> , \RAM<0><4> ,
         \RAM<0><3> , \RAM<0><2> , \RAM<0><1> , \RAM<0><0> , n66, n3519, n3520,
         n3521, n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530,
         n3531, n3532, n3533, n3534, n3535, n3536, n3538, n3539, n3540, n3541,
         n3542, n3543, n3544, n3545, n3546, n3548, n3549, n3550, n3551, n3552,
         n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3562, n3563, n3564,
         n3567, n3568, n3570, n3571, n3572, n3573, n3574, n3575, n3577, n3578,
         n3579, n3580, n3581, n3565, n3569, n3582, n3583, n3560, n3561, n3566,
         n3576, n2056, n2057, n2058, n2059, n2060, n2061, n2063, n2064, n2065,
         n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075,
         n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085,
         n2086, n2087, n2088, n2090, n2091, n2092, n2093, n2094, n2095, n2096,
         n2097, n2098, n2099, n2101, n2102, n2103, n2104, n2105, n2106, n2107,
         n2108, n2109, n2110, n2112, n2113, n2114, n2115, n2116, n2117, n2118,
         n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128,
         n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138,
         n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148,
         n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158,
         n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168,
         n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178,
         n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188,
         n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198,
         n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208,
         n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218,
         n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228,
         n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238,
         n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248,
         n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258,
         n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268,
         n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278,
         n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288,
         n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298,
         n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308,
         n2309, n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318,
         n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328,
         n2329, n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338,
         n2339, n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348,
         n2349, n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358,
         n2359, n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368,
         n2369, n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378,
         n2379, n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388,
         n2389, n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398,
         n2399, n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408,
         n2409, n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418,
         n2419, n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428,
         n2429, n2430, n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438,
         n2439, n2440, n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448,
         n2449, n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458,
         n2459, n2460, n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468,
         n2469, n2470, n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478,
         n2479, n2480, n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488,
         n2489, n2490, n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498,
         n2499, n2500, n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508,
         n2509, n2510, n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518,
         n2519, n2520, n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528,
         n2529, n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538,
         n2539, n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548,
         n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558,
         n2559, n2560, n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568,
         n2569, n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578,
         n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588,
         n2589, n2590, n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598,
         n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608,
         n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618,
         n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628,
         n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638,
         n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648,
         n2649, n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658,
         n2659, n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668,
         n2669, n2670, n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678,
         n2679, n2680, n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2688,
         n2689, n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698,
         n2699, n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2708,
         n2709, n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718,
         n2719, n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728,
         n2729, n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737, n2738,
         n2739, n2740, n2741, n2742, n2743, n2744, n2745, n2746, n2747, n2748,
         n2749, n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758,
         n2759, n2760, n2761, n2762, n2763, n2764, n2765, n2766, n2767, n2768,
         n2769, n2770, n2771, n2772, n2773, n2774, n2775, n2776, n2777, n2778,
         n2779, n2780, n2781, n2782, n2783, n2784, n2785, n2786, n2787, n2788,
         n2789, n2790, n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798,
         n2799, n2800, n2801, n2802, n2803, n2804, n2805, n2806, n2807, n2808,
         n2809, n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817, n2818,
         n2819, n2820, n2821, n2822, n2823, n2824, n2825, n2826, n2827, n2828,
         n2829, n2830, n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2838,
         n2839, n2840, n2841, n2842, n2843, n2844, n2845, n2846, n2847, n2848,
         n2849, n2850, n2851, n2852, n2853, n2854, n2855, n2856, n2857, n2858,
         n2859, n2860, n2861, n2862, n2863, n2864, n2865, n2866, n2867, n2868,
         n2869, n2870, n2871, n2872, n2873, n2874, n2875, n2876, n2877, n2878,
         n2879, n2880, n2881, n2882, n2883, n2884, n2885, n2886, n2887, n2888,
         n2889, n2890, n2891, n2892, n2893, n2894, n2895, n2896, n2897, n2898,
         n2899, n2900, n2901, n2902, n2903, n2904, n2905, n2906, n2907, n2908,
         n2909, n2910, n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2918,
         n2919, n2920, n2921, n2922, n2923, n2924, n2925, n2926, n2927, n2928,
         n2929, n2930, n2931, n2932, n2933, n2934, n2935, n2936, n2937, n2938,
         n2939, n2940, n2941, n2942, n2943, n2944, n2945, n2946, n2947, n2948,
         n2949, n2950, n2951, n2952, n2953, n2954, n2955, n2956, n2957, n2958,
         n2959, n2960, n2961, n2962, n2963, n2964, n2965, n2966, n2967, n2968,
         n2969, n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977, n2978,
         n2979, n2980, n2981, n2982, n2983, n2984, n2985, n2986, n2987, n2988,
         n2989, n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998,
         n2999, n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007, n3008,
         n3009, n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017, n3018,
         n3019, n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027, n3028,
         n3029, n3030, n3031, n3032, n3033, n3034, n3035, n3036, n3037, n3038,
         n3039, n3040, n3041, n3042, n3043, n3044, n3045, n3046, n3047, n3048,
         n3049, n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057, n3058,
         n3059, n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067, n3068,
         n3069, n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078,
         n3079, n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3088,
         n3089, n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097, n3098,
         n3099, n3100, n3101, n3102, n3103, n3104, n3105, n3106, n3107, n3108,
         n3109, n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118,
         n3119, n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3127, n3128,
         n3129, n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3138,
         n3139, n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147, n3148,
         n3149, n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157, n3158,
         n3159, n3160, n3161, n3162, n3163, n3164, n3165, n3166, n3167, n3168,
         n3169, n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178,
         n3179, n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188,
         n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198,
         n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208,
         n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218,
         n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228,
         n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238,
         n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248,
         n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258,
         n3259, n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268,
         n3269, n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278,
         n3279, n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288,
         n3289, n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298,
         n3299, n3300, n3301, n3302, n3303, n3304, n3305, n3306, n3307, n3308,
         n3309, n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318,
         n3319, n3320, n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328,
         n3329, n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338,
         n3339, n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348,
         n3349, n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358,
         n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368,
         n3369, n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378,
         n3379, n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388,
         n3389, n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398,
         n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408,
         n3409, n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418,
         n3419, n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428,
         n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438,
         n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448,
         n3449, n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458,
         n3459, n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468,
         n3469, n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478,
         n3479, n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487, n3488,
         n3489, n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497, n3498,
         n3499, n3500, n3501, n3502, n3503, n3504, n3505, n3506, n3507, n3508,
         n3509, n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518,
         n3537, n3547, n16074, n16075, n16076, n16077, n18126, n18127, n18128,
         n18129, n18130, n18131, n18132, n18133, n18134, n18135, n18136,
         n18137, n18138, n18139, n18140, n18141, n18142, n18143, n18144,
         n18145, n18146, n18147, n18148, n18149, n18150, n18151, n18152,
         n18153, n18154, n18155, n18156, n18157, n18158, n18159, n18160,
         n18161, n18162, n18163, n18164, n18165, n18166, n18167, n18168,
         n18169, n18170, n18171, n18172, n18173, n18174, n18175, n18176,
         n18177, n18178, n18179, n18180, n18181, n18182, n18183, n18184,
         n18185, n18186, n18187, n18188, n18189, n18190, n18191, n18192,
         n18193, n18194, n18195, n18196, n18197, n18198, n18199, n18200,
         n18201, n18202, n18203, n18204, n18205, n18206, n18207, n18208,
         n18209, n18210, n18211, n18212, n18213, n18214, n18215, n18216,
         n18217, n18218, n18219, n18220, n18221, n18222, n18223, n18224,
         n18225, n18226, n18227, n18228, n18229, n18230, n18231, n18232,
         n18233, n18234, n18235, n18236, n18237, n18238, n18239, n18240,
         n18241, n18242, n18243, n18244, n18245, n18246, n18247, n18248,
         n18249, n18250, n18251, n18252, n18253, n18254, n18255, n18256,
         n18257, n18258, n18259, n18260, n18261, n18262, n18263, n18264,
         n18265, n18266, n18267, n18268, n18269, n18270, n18271, n18272,
         n18273, n18274, n18275, n18276, n18277, n18278, n18279, n18280,
         n18281, n18282, n18283, n18284, n18285, n18286, n18287, n18288,
         n18289, n18290, n18291, n18292, n18293, n18294, n18295, n18296,
         n18297, n18298, n18299, n18300, n18301, n18302, n18303, n18304,
         n18305, n18306, n18307, n18308, n18309, n18310, n18311, n18312,
         n18313, n18314, n18315, n18316, n18317, n18318, n18319, n18320,
         n18321, n18322, n18323, n18324, n18325, n18326, n18327, n18328,
         n18329, n18330, n18331, n18332, n18333, n18334, n18335, n18336,
         n18337, n18338, n18339, n18340, n18341, n18342, n18343, n18344,
         n18345, n18346, n18347, n18348, n18349, n18350, n18351, n18352,
         n18353, n18354, n18355, n18356, n18357, n18358, n18359, n18360,
         n18361, n18362, n18363, n18364, n18365, n18366, n18367, n18368,
         n18369, n18370, n18371, n18372, n18373, n18374, n18375, n18376,
         n18377, n18378, n18379, n18380, n18381, n18382, n18383, n18384,
         n18385, n18386, n18387, n18388, n18389, n18390, n18391, n18392,
         n18393, n18394, n18395, n18396, n18397, n18398, n18399, n18400,
         n18401, n18402, n18403, n18404, n18405, n18406, n18407, n18408,
         n18409, n18410, n18411, n18412, n18413, n18414, n18415, n18416,
         n18417, n18418, n18419, n18420, n18421, n18422, n18423, n18424,
         n18425, n18426, n18427, n18428, n18429, n18430, n18431, n18432,
         n18433, n18434, n18435, n18436, n18437, n18438, n18439, n18440,
         n18441, n18442, n18443, n18444, n18445, n18446, n18447, n18448,
         n18449, n18450, n18451, n18452, n18453, n18454, n18455, n18456,
         n18457, n18458, n18459, n18460, n18461, n18462, n18463, n18464,
         n18465, n18466, n18467, n18468, n18469, n18470, n18471, n18472,
         n18473, n18474, n18475, n18476, n18477, n18478, n18479, n18480,
         n18481, n18482, n18483, n18484, n18485, n18486, n18487, n18488,
         n18489, n18490, n18491, n18492, n18493, n18494, n18495, n18496,
         n18497, n18498, n18499, n18500, n18501, n18502, n18503, n18504,
         n18505, n18506, n18507, n18508, n18509, n18510, n18511, n18512,
         n18513, n18514, n18515, n18516, n18517, n18518, n18519, n18520,
         n18521, n18522, n18523, n18524, n18525, n18526, n18527, n18528,
         n18529, n18530, n18531, n18532, n18533, n18534, n18535, n18536,
         n18537, n18538, n18539, n18540, n18541, n18542, n18543, n18544,
         n18545, n18546, n18547, n18548, n18549, n18550, n18551, n18552,
         n18553, n18554, n18555, n18556, n18557, n18558, n18559, n18560,
         n18561, n18562, n18563, n18564, n18565, n18566, n18567, n18568,
         n18569, n18570, n18571;
  assign N32 = \a<2> ;
  assign N33 = \a<3> ;
  assign N34 = \a<4> ;
  assign N35 = \a<5> ;
  assign N36 = \a<6> ;
  assign N37 = \a<7> ;

  EDFFX1 \RAM_reg<57><31>  ( .D(n18564), .E(n18327), .CK(clk), .Q(
        \RAM<57><31> ) );
  EDFFX1 \RAM_reg<57><30>  ( .D(n18560), .E(n18327), .CK(clk), .Q(
        \RAM<57><30> ) );
  EDFFX1 \RAM_reg<57><29>  ( .D(n18556), .E(n18327), .CK(clk), .Q(
        \RAM<57><29> ) );
  EDFFX1 \RAM_reg<57><28>  ( .D(n18552), .E(n18327), .CK(clk), .Q(
        \RAM<57><28> ) );
  EDFFX1 \RAM_reg<57><27>  ( .D(n18548), .E(n18327), .CK(clk), .Q(
        \RAM<57><27> ) );
  EDFFX1 \RAM_reg<57><26>  ( .D(n18544), .E(n18327), .CK(clk), .Q(
        \RAM<57><26> ) );
  EDFFX1 \RAM_reg<57><25>  ( .D(n18540), .E(n18327), .CK(clk), .Q(
        \RAM<57><25> ) );
  EDFFX1 \RAM_reg<57><24>  ( .D(n18536), .E(n18327), .CK(clk), .Q(
        \RAM<57><24> ) );
  EDFFX1 \RAM_reg<57><23>  ( .D(n18532), .E(n18327), .CK(clk), .Q(
        \RAM<57><23> ) );
  EDFFX1 \RAM_reg<57><22>  ( .D(n18528), .E(n18327), .CK(clk), .Q(
        \RAM<57><22> ) );
  EDFFX1 \RAM_reg<57><21>  ( .D(n18524), .E(n18327), .CK(clk), .Q(
        \RAM<57><21> ) );
  EDFFX1 \RAM_reg<57><20>  ( .D(n18520), .E(n18327), .CK(clk), .Q(
        \RAM<57><20> ) );
  EDFFX1 \RAM_reg<57><19>  ( .D(n18516), .E(n18328), .CK(clk), .Q(
        \RAM<57><19> ) );
  EDFFX1 \RAM_reg<57><18>  ( .D(n18512), .E(n18328), .CK(clk), .Q(
        \RAM<57><18> ) );
  EDFFX1 \RAM_reg<57><17>  ( .D(n18508), .E(n18328), .CK(clk), .Q(
        \RAM<57><17> ) );
  EDFFX1 \RAM_reg<57><16>  ( .D(n18504), .E(n18328), .CK(clk), .Q(
        \RAM<57><16> ) );
  EDFFX1 \RAM_reg<57><15>  ( .D(n18500), .E(n18328), .CK(clk), .Q(
        \RAM<57><15> ) );
  EDFFX1 \RAM_reg<57><14>  ( .D(n18496), .E(n18328), .CK(clk), .Q(
        \RAM<57><14> ) );
  EDFFX1 \RAM_reg<57><13>  ( .D(n18492), .E(n18328), .CK(clk), .Q(
        \RAM<57><13> ) );
  EDFFX1 \RAM_reg<57><12>  ( .D(n18488), .E(n18328), .CK(clk), .Q(
        \RAM<57><12> ) );
  EDFFX1 \RAM_reg<57><11>  ( .D(n18484), .E(n18328), .CK(clk), .Q(
        \RAM<57><11> ) );
  EDFFX1 \RAM_reg<57><10>  ( .D(n18480), .E(n18328), .CK(clk), .Q(
        \RAM<57><10> ) );
  EDFFX1 \RAM_reg<57><9>  ( .D(n18476), .E(n18328), .CK(clk), .Q(\RAM<57><9> )
         );
  EDFFX1 \RAM_reg<57><8>  ( .D(n18472), .E(n18328), .CK(clk), .Q(\RAM<57><8> )
         );
  EDFFX1 \RAM_reg<57><7>  ( .D(n18468), .E(n3556), .CK(clk), .Q(\RAM<57><7> )
         );
  EDFFX1 \RAM_reg<57><6>  ( .D(n18464), .E(n3556), .CK(clk), .Q(\RAM<57><6> )
         );
  EDFFX1 \RAM_reg<57><5>  ( .D(n18460), .E(n18327), .CK(clk), .Q(\RAM<57><5> )
         );
  EDFFX1 \RAM_reg<57><4>  ( .D(n18456), .E(n18328), .CK(clk), .Q(\RAM<57><4> )
         );
  EDFFX1 \RAM_reg<57><3>  ( .D(n18452), .E(n18327), .CK(clk), .Q(\RAM<57><3> )
         );
  EDFFX1 \RAM_reg<57><2>  ( .D(n18448), .E(n18328), .CK(clk), .Q(\RAM<57><2> )
         );
  EDFFX1 \RAM_reg<57><1>  ( .D(n18444), .E(n18327), .CK(clk), .Q(\RAM<57><1> )
         );
  EDFFX1 \RAM_reg<57><0>  ( .D(n18440), .E(n18328), .CK(clk), .Q(\RAM<57><0> )
         );
  EDFFX1 \RAM_reg<49><31>  ( .D(n18562), .E(n18390), .CK(clk), .Q(
        \RAM<49><31> ) );
  EDFFX1 \RAM_reg<49><30>  ( .D(n18558), .E(n18390), .CK(clk), .Q(
        \RAM<49><30> ) );
  EDFFX1 \RAM_reg<49><29>  ( .D(n18554), .E(n18390), .CK(clk), .Q(
        \RAM<49><29> ) );
  EDFFX1 \RAM_reg<49><28>  ( .D(n18550), .E(n18390), .CK(clk), .Q(
        \RAM<49><28> ) );
  EDFFX1 \RAM_reg<49><27>  ( .D(n18546), .E(n18390), .CK(clk), .Q(
        \RAM<49><27> ) );
  EDFFX1 \RAM_reg<49><26>  ( .D(n18542), .E(n18390), .CK(clk), .Q(
        \RAM<49><26> ) );
  EDFFX1 \RAM_reg<49><25>  ( .D(n18538), .E(n18390), .CK(clk), .Q(
        \RAM<49><25> ) );
  EDFFX1 \RAM_reg<49><24>  ( .D(n18534), .E(n18390), .CK(clk), .Q(
        \RAM<49><24> ) );
  EDFFX1 \RAM_reg<49><23>  ( .D(n18530), .E(n18390), .CK(clk), .Q(
        \RAM<49><23> ) );
  EDFFX1 \RAM_reg<49><22>  ( .D(n18526), .E(n18390), .CK(clk), .Q(
        \RAM<49><22> ) );
  EDFFX1 \RAM_reg<49><21>  ( .D(n18522), .E(n18390), .CK(clk), .Q(
        \RAM<49><21> ) );
  EDFFX1 \RAM_reg<49><20>  ( .D(n18518), .E(n18390), .CK(clk), .Q(
        \RAM<49><20> ) );
  EDFFX1 \RAM_reg<49><19>  ( .D(n18514), .E(n18391), .CK(clk), .Q(
        \RAM<49><19> ) );
  EDFFX1 \RAM_reg<49><18>  ( .D(n18510), .E(n18391), .CK(clk), .Q(
        \RAM<49><18> ) );
  EDFFX1 \RAM_reg<49><17>  ( .D(n18506), .E(n18391), .CK(clk), .Q(
        \RAM<49><17> ) );
  EDFFX1 \RAM_reg<49><16>  ( .D(n18502), .E(n18391), .CK(clk), .Q(
        \RAM<49><16> ) );
  EDFFX1 \RAM_reg<49><15>  ( .D(n18498), .E(n18391), .CK(clk), .Q(
        \RAM<49><15> ) );
  EDFFX1 \RAM_reg<49><14>  ( .D(n18494), .E(n18391), .CK(clk), .Q(
        \RAM<49><14> ) );
  EDFFX1 \RAM_reg<49><13>  ( .D(n18490), .E(n18391), .CK(clk), .Q(
        \RAM<49><13> ) );
  EDFFX1 \RAM_reg<49><12>  ( .D(n18486), .E(n18391), .CK(clk), .Q(
        \RAM<49><12> ) );
  EDFFX1 \RAM_reg<49><11>  ( .D(n18482), .E(n18391), .CK(clk), .Q(
        \RAM<49><11> ) );
  EDFFX1 \RAM_reg<49><10>  ( .D(n18478), .E(n18391), .CK(clk), .Q(
        \RAM<49><10> ) );
  EDFFX1 \RAM_reg<49><9>  ( .D(n18474), .E(n18391), .CK(clk), .Q(\RAM<49><9> )
         );
  EDFFX1 \RAM_reg<49><8>  ( .D(n18470), .E(n18391), .CK(clk), .Q(\RAM<49><8> )
         );
  EDFFX1 \RAM_reg<49><7>  ( .D(n18466), .E(n3533), .CK(clk), .Q(\RAM<49><7> )
         );
  EDFFX1 \RAM_reg<49><6>  ( .D(n18462), .E(n3533), .CK(clk), .Q(\RAM<49><6> )
         );
  EDFFX1 \RAM_reg<49><5>  ( .D(n18458), .E(n18390), .CK(clk), .Q(\RAM<49><5> )
         );
  EDFFX1 \RAM_reg<49><4>  ( .D(n18454), .E(n18391), .CK(clk), .Q(\RAM<49><4> )
         );
  EDFFX1 \RAM_reg<49><3>  ( .D(n18450), .E(n18390), .CK(clk), .Q(\RAM<49><3> )
         );
  EDFFX1 \RAM_reg<49><2>  ( .D(n18446), .E(n18391), .CK(clk), .Q(\RAM<49><2> )
         );
  EDFFX1 \RAM_reg<49><1>  ( .D(n18442), .E(n18390), .CK(clk), .Q(\RAM<49><1> )
         );
  EDFFX1 \RAM_reg<49><0>  ( .D(n18438), .E(n18391), .CK(clk), .Q(\RAM<49><0> )
         );
  EDFFX1 \RAM_reg<41><31>  ( .D(n18563), .E(n18384), .CK(clk), .Q(
        \RAM<41><31> ) );
  EDFFX1 \RAM_reg<41><30>  ( .D(n18559), .E(n18384), .CK(clk), .Q(
        \RAM<41><30> ) );
  EDFFX1 \RAM_reg<41><29>  ( .D(n18555), .E(n18384), .CK(clk), .Q(
        \RAM<41><29> ) );
  EDFFX1 \RAM_reg<41><28>  ( .D(n18551), .E(n18384), .CK(clk), .Q(
        \RAM<41><28> ) );
  EDFFX1 \RAM_reg<41><27>  ( .D(n18547), .E(n18384), .CK(clk), .Q(
        \RAM<41><27> ) );
  EDFFX1 \RAM_reg<41><26>  ( .D(n18543), .E(n18384), .CK(clk), .Q(
        \RAM<41><26> ) );
  EDFFX1 \RAM_reg<41><25>  ( .D(n18539), .E(n18384), .CK(clk), .Q(
        \RAM<41><25> ) );
  EDFFX1 \RAM_reg<41><24>  ( .D(n18535), .E(n18384), .CK(clk), .Q(
        \RAM<41><24> ) );
  EDFFX1 \RAM_reg<41><23>  ( .D(n18531), .E(n18384), .CK(clk), .Q(
        \RAM<41><23> ) );
  EDFFX1 \RAM_reg<41><22>  ( .D(n18527), .E(n18384), .CK(clk), .Q(
        \RAM<41><22> ) );
  EDFFX1 \RAM_reg<41><21>  ( .D(n18523), .E(n18384), .CK(clk), .Q(
        \RAM<41><21> ) );
  EDFFX1 \RAM_reg<41><20>  ( .D(n18519), .E(n18384), .CK(clk), .Q(
        \RAM<41><20> ) );
  EDFFX1 \RAM_reg<41><19>  ( .D(n18515), .E(n18385), .CK(clk), .Q(
        \RAM<41><19> ) );
  EDFFX1 \RAM_reg<41><18>  ( .D(n18511), .E(n18385), .CK(clk), .Q(
        \RAM<41><18> ) );
  EDFFX1 \RAM_reg<41><17>  ( .D(n18507), .E(n18385), .CK(clk), .Q(
        \RAM<41><17> ) );
  EDFFX1 \RAM_reg<41><16>  ( .D(n18503), .E(n18385), .CK(clk), .Q(
        \RAM<41><16> ) );
  EDFFX1 \RAM_reg<41><15>  ( .D(n18499), .E(n18385), .CK(clk), .Q(
        \RAM<41><15> ) );
  EDFFX1 \RAM_reg<41><14>  ( .D(n18495), .E(n18385), .CK(clk), .Q(
        \RAM<41><14> ) );
  EDFFX1 \RAM_reg<41><13>  ( .D(n18491), .E(n18385), .CK(clk), .Q(
        \RAM<41><13> ) );
  EDFFX1 \RAM_reg<41><12>  ( .D(n18487), .E(n18385), .CK(clk), .Q(
        \RAM<41><12> ) );
  EDFFX1 \RAM_reg<41><11>  ( .D(n18483), .E(n18385), .CK(clk), .Q(
        \RAM<41><11> ) );
  EDFFX1 \RAM_reg<41><10>  ( .D(n18479), .E(n18385), .CK(clk), .Q(
        \RAM<41><10> ) );
  EDFFX1 \RAM_reg<41><9>  ( .D(n18475), .E(n18385), .CK(clk), .Q(\RAM<41><9> )
         );
  EDFFX1 \RAM_reg<41><8>  ( .D(n18471), .E(n18385), .CK(clk), .Q(\RAM<41><8> )
         );
  EDFFX1 \RAM_reg<41><7>  ( .D(n18467), .E(n3535), .CK(clk), .Q(\RAM<41><7> )
         );
  EDFFX1 \RAM_reg<41><6>  ( .D(n18463), .E(n3535), .CK(clk), .Q(\RAM<41><6> )
         );
  EDFFX1 \RAM_reg<41><5>  ( .D(n18459), .E(n18384), .CK(clk), .Q(\RAM<41><5> )
         );
  EDFFX1 \RAM_reg<41><4>  ( .D(n18455), .E(n18385), .CK(clk), .Q(\RAM<41><4> )
         );
  EDFFX1 \RAM_reg<41><3>  ( .D(n18451), .E(n18384), .CK(clk), .Q(\RAM<41><3> )
         );
  EDFFX1 \RAM_reg<41><2>  ( .D(n18447), .E(n18385), .CK(clk), .Q(\RAM<41><2> )
         );
  EDFFX1 \RAM_reg<41><1>  ( .D(n18443), .E(n18384), .CK(clk), .Q(\RAM<41><1> )
         );
  EDFFX1 \RAM_reg<41><0>  ( .D(n18439), .E(n18385), .CK(clk), .Q(\RAM<41><0> )
         );
  EDFFX1 \RAM_reg<33><31>  ( .D(\wd<31> ), .E(n18339), .CK(clk), .Q(
        \RAM<33><31> ) );
  EDFFX1 \RAM_reg<33><30>  ( .D(\wd<30> ), .E(n18339), .CK(clk), .Q(
        \RAM<33><30> ) );
  EDFFX1 \RAM_reg<33><29>  ( .D(\wd<29> ), .E(n18339), .CK(clk), .Q(
        \RAM<33><29> ) );
  EDFFX1 \RAM_reg<33><28>  ( .D(\wd<28> ), .E(n18339), .CK(clk), .Q(
        \RAM<33><28> ) );
  EDFFX1 \RAM_reg<33><27>  ( .D(\wd<27> ), .E(n18339), .CK(clk), .Q(
        \RAM<33><27> ) );
  EDFFX1 \RAM_reg<33><26>  ( .D(\wd<26> ), .E(n18339), .CK(clk), .Q(
        \RAM<33><26> ) );
  EDFFX1 \RAM_reg<33><25>  ( .D(\wd<25> ), .E(n18339), .CK(clk), .Q(
        \RAM<33><25> ) );
  EDFFX1 \RAM_reg<33><24>  ( .D(\wd<24> ), .E(n18339), .CK(clk), .Q(
        \RAM<33><24> ) );
  EDFFX1 \RAM_reg<33><23>  ( .D(\wd<23> ), .E(n18339), .CK(clk), .Q(
        \RAM<33><23> ) );
  EDFFX1 \RAM_reg<33><22>  ( .D(\wd<22> ), .E(n18339), .CK(clk), .Q(
        \RAM<33><22> ) );
  EDFFX1 \RAM_reg<33><21>  ( .D(\wd<21> ), .E(n18339), .CK(clk), .Q(
        \RAM<33><21> ) );
  EDFFX1 \RAM_reg<33><20>  ( .D(\wd<20> ), .E(n18339), .CK(clk), .Q(
        \RAM<33><20> ) );
  EDFFX1 \RAM_reg<33><19>  ( .D(\wd<19> ), .E(n18340), .CK(clk), .Q(
        \RAM<33><19> ) );
  EDFFX1 \RAM_reg<33><18>  ( .D(\wd<18> ), .E(n18340), .CK(clk), .Q(
        \RAM<33><18> ) );
  EDFFX1 \RAM_reg<33><17>  ( .D(\wd<17> ), .E(n18340), .CK(clk), .Q(
        \RAM<33><17> ) );
  EDFFX1 \RAM_reg<33><16>  ( .D(\wd<16> ), .E(n18340), .CK(clk), .Q(
        \RAM<33><16> ) );
  EDFFX1 \RAM_reg<33><15>  ( .D(\wd<15> ), .E(n18340), .CK(clk), .Q(
        \RAM<33><15> ) );
  EDFFX1 \RAM_reg<33><14>  ( .D(\wd<14> ), .E(n18340), .CK(clk), .Q(
        \RAM<33><14> ) );
  EDFFX1 \RAM_reg<33><13>  ( .D(\wd<13> ), .E(n18340), .CK(clk), .Q(
        \RAM<33><13> ) );
  EDFFX1 \RAM_reg<33><12>  ( .D(\wd<12> ), .E(n18340), .CK(clk), .Q(
        \RAM<33><12> ) );
  EDFFX1 \RAM_reg<33><11>  ( .D(\wd<11> ), .E(n18340), .CK(clk), .Q(
        \RAM<33><11> ) );
  EDFFX1 \RAM_reg<33><10>  ( .D(\wd<10> ), .E(n18340), .CK(clk), .Q(
        \RAM<33><10> ) );
  EDFFX1 \RAM_reg<33><9>  ( .D(\wd<9> ), .E(n18340), .CK(clk), .Q(\RAM<33><9> ) );
  EDFFX1 \RAM_reg<33><8>  ( .D(\wd<8> ), .E(n18340), .CK(clk), .Q(\RAM<33><8> ) );
  EDFFX1 \RAM_reg<33><7>  ( .D(\wd<7> ), .E(n3552), .CK(clk), .Q(\RAM<33><7> )
         );
  EDFFX1 \RAM_reg<33><6>  ( .D(\wd<6> ), .E(n3552), .CK(clk), .Q(\RAM<33><6> )
         );
  EDFFX1 \RAM_reg<33><5>  ( .D(\wd<5> ), .E(n18339), .CK(clk), .Q(\RAM<33><5> ) );
  EDFFX1 \RAM_reg<33><4>  ( .D(\wd<4> ), .E(n18340), .CK(clk), .Q(\RAM<33><4> ) );
  EDFFX1 \RAM_reg<33><3>  ( .D(\wd<3> ), .E(n18339), .CK(clk), .Q(\RAM<33><3> ) );
  EDFFX1 \RAM_reg<33><2>  ( .D(\wd<2> ), .E(n18340), .CK(clk), .Q(\RAM<33><2> ) );
  EDFFX1 \RAM_reg<33><1>  ( .D(\wd<1> ), .E(n18339), .CK(clk), .Q(\RAM<33><1> ) );
  EDFFX1 \RAM_reg<33><0>  ( .D(\wd<0> ), .E(n18340), .CK(clk), .Q(\RAM<33><0> ) );
  EDFFX1 \RAM_reg<25><31>  ( .D(n18562), .E(n18426), .CK(clk), .Q(
        \RAM<25><31> ) );
  EDFFX1 \RAM_reg<25><30>  ( .D(n18558), .E(n18426), .CK(clk), .Q(
        \RAM<25><30> ) );
  EDFFX1 \RAM_reg<25><29>  ( .D(n18554), .E(n18426), .CK(clk), .Q(
        \RAM<25><29> ) );
  EDFFX1 \RAM_reg<25><28>  ( .D(n18550), .E(n18426), .CK(clk), .Q(
        \RAM<25><28> ) );
  EDFFX1 \RAM_reg<25><27>  ( .D(n18546), .E(n18426), .CK(clk), .Q(
        \RAM<25><27> ) );
  EDFFX1 \RAM_reg<25><26>  ( .D(n18542), .E(n18426), .CK(clk), .Q(
        \RAM<25><26> ) );
  EDFFX1 \RAM_reg<25><25>  ( .D(n18538), .E(n18426), .CK(clk), .Q(
        \RAM<25><25> ) );
  EDFFX1 \RAM_reg<25><24>  ( .D(n18534), .E(n18426), .CK(clk), .Q(
        \RAM<25><24> ) );
  EDFFX1 \RAM_reg<25><23>  ( .D(n18530), .E(n18426), .CK(clk), .Q(
        \RAM<25><23> ) );
  EDFFX1 \RAM_reg<25><22>  ( .D(n18526), .E(n18426), .CK(clk), .Q(
        \RAM<25><22> ) );
  EDFFX1 \RAM_reg<25><21>  ( .D(n18522), .E(n18426), .CK(clk), .Q(
        \RAM<25><21> ) );
  EDFFX1 \RAM_reg<25><20>  ( .D(n18518), .E(n18426), .CK(clk), .Q(
        \RAM<25><20> ) );
  EDFFX1 \RAM_reg<25><19>  ( .D(n18514), .E(n18427), .CK(clk), .Q(
        \RAM<25><19> ) );
  EDFFX1 \RAM_reg<25><18>  ( .D(n18510), .E(n18427), .CK(clk), .Q(
        \RAM<25><18> ) );
  EDFFX1 \RAM_reg<25><17>  ( .D(n18506), .E(n18427), .CK(clk), .Q(
        \RAM<25><17> ) );
  EDFFX1 \RAM_reg<25><16>  ( .D(n18502), .E(n18427), .CK(clk), .Q(
        \RAM<25><16> ) );
  EDFFX1 \RAM_reg<25><15>  ( .D(n18498), .E(n18427), .CK(clk), .Q(
        \RAM<25><15> ) );
  EDFFX1 \RAM_reg<25><14>  ( .D(n18494), .E(n18427), .CK(clk), .Q(
        \RAM<25><14> ) );
  EDFFX1 \RAM_reg<25><13>  ( .D(n18490), .E(n18427), .CK(clk), .Q(
        \RAM<25><13> ) );
  EDFFX1 \RAM_reg<25><12>  ( .D(n18486), .E(n18427), .CK(clk), .Q(
        \RAM<25><12> ) );
  EDFFX1 \RAM_reg<25><11>  ( .D(n18482), .E(n18427), .CK(clk), .Q(
        \RAM<25><11> ) );
  EDFFX1 \RAM_reg<25><10>  ( .D(n18478), .E(n18427), .CK(clk), .Q(
        \RAM<25><10> ) );
  EDFFX1 \RAM_reg<25><9>  ( .D(n18474), .E(n18427), .CK(clk), .Q(\RAM<25><9> )
         );
  EDFFX1 \RAM_reg<25><8>  ( .D(n18470), .E(n18427), .CK(clk), .Q(\RAM<25><8> )
         );
  EDFFX1 \RAM_reg<25><7>  ( .D(n18466), .E(n3521), .CK(clk), .Q(\RAM<25><7> )
         );
  EDFFX1 \RAM_reg<25><6>  ( .D(n18462), .E(n3521), .CK(clk), .Q(\RAM<25><6> )
         );
  EDFFX1 \RAM_reg<25><5>  ( .D(n18458), .E(n18426), .CK(clk), .Q(\RAM<25><5> )
         );
  EDFFX1 \RAM_reg<25><4>  ( .D(n18454), .E(n18427), .CK(clk), .Q(\RAM<25><4> )
         );
  EDFFX1 \RAM_reg<25><3>  ( .D(n18450), .E(n18426), .CK(clk), .Q(\RAM<25><3> )
         );
  EDFFX1 \RAM_reg<25><2>  ( .D(n18446), .E(n18427), .CK(clk), .Q(\RAM<25><2> )
         );
  EDFFX1 \RAM_reg<25><1>  ( .D(n18442), .E(n18426), .CK(clk), .Q(\RAM<25><1> )
         );
  EDFFX1 \RAM_reg<25><0>  ( .D(n18438), .E(n18427), .CK(clk), .Q(\RAM<25><0> )
         );
  EDFFX1 \RAM_reg<17><31>  ( .D(n18563), .E(n18372), .CK(clk), .Q(
        \RAM<17><31> ) );
  EDFFX1 \RAM_reg<17><30>  ( .D(n18559), .E(n18372), .CK(clk), .Q(
        \RAM<17><30> ) );
  EDFFX1 \RAM_reg<17><29>  ( .D(n18555), .E(n18372), .CK(clk), .Q(
        \RAM<17><29> ) );
  EDFFX1 \RAM_reg<17><28>  ( .D(n18551), .E(n18372), .CK(clk), .Q(
        \RAM<17><28> ) );
  EDFFX1 \RAM_reg<17><27>  ( .D(n18547), .E(n18372), .CK(clk), .Q(
        \RAM<17><27> ) );
  EDFFX1 \RAM_reg<17><26>  ( .D(n18543), .E(n18372), .CK(clk), .Q(
        \RAM<17><26> ) );
  EDFFX1 \RAM_reg<17><25>  ( .D(n18539), .E(n18372), .CK(clk), .Q(
        \RAM<17><25> ) );
  EDFFX1 \RAM_reg<17><24>  ( .D(n18535), .E(n18372), .CK(clk), .Q(
        \RAM<17><24> ) );
  EDFFX1 \RAM_reg<17><23>  ( .D(n18531), .E(n18372), .CK(clk), .Q(
        \RAM<17><23> ) );
  EDFFX1 \RAM_reg<17><22>  ( .D(n18527), .E(n18372), .CK(clk), .Q(
        \RAM<17><22> ) );
  EDFFX1 \RAM_reg<17><21>  ( .D(n18523), .E(n18372), .CK(clk), .Q(
        \RAM<17><21> ) );
  EDFFX1 \RAM_reg<17><20>  ( .D(n18519), .E(n18372), .CK(clk), .Q(
        \RAM<17><20> ) );
  EDFFX1 \RAM_reg<17><19>  ( .D(n18515), .E(n18373), .CK(clk), .Q(
        \RAM<17><19> ) );
  EDFFX1 \RAM_reg<17><18>  ( .D(n18511), .E(n18373), .CK(clk), .Q(
        \RAM<17><18> ) );
  EDFFX1 \RAM_reg<17><17>  ( .D(n18507), .E(n18373), .CK(clk), .Q(
        \RAM<17><17> ) );
  EDFFX1 \RAM_reg<17><16>  ( .D(n18503), .E(n18373), .CK(clk), .Q(
        \RAM<17><16> ) );
  EDFFX1 \RAM_reg<17><15>  ( .D(n18499), .E(n18373), .CK(clk), .Q(
        \RAM<17><15> ) );
  EDFFX1 \RAM_reg<17><14>  ( .D(n18495), .E(n18373), .CK(clk), .Q(
        \RAM<17><14> ) );
  EDFFX1 \RAM_reg<17><13>  ( .D(n18491), .E(n18373), .CK(clk), .Q(
        \RAM<17><13> ) );
  EDFFX1 \RAM_reg<17><12>  ( .D(n18487), .E(n18373), .CK(clk), .Q(
        \RAM<17><12> ) );
  EDFFX1 \RAM_reg<17><11>  ( .D(n18483), .E(n18373), .CK(clk), .Q(
        \RAM<17><11> ) );
  EDFFX1 \RAM_reg<17><10>  ( .D(n18479), .E(n18373), .CK(clk), .Q(
        \RAM<17><10> ) );
  EDFFX1 \RAM_reg<17><9>  ( .D(n18475), .E(n18373), .CK(clk), .Q(\RAM<17><9> )
         );
  EDFFX1 \RAM_reg<17><8>  ( .D(n18471), .E(n18373), .CK(clk), .Q(\RAM<17><8> )
         );
  EDFFX1 \RAM_reg<17><7>  ( .D(n18467), .E(n3540), .CK(clk), .Q(\RAM<17><7> )
         );
  EDFFX1 \RAM_reg<17><6>  ( .D(n18463), .E(n3540), .CK(clk), .Q(\RAM<17><6> )
         );
  EDFFX1 \RAM_reg<17><5>  ( .D(n18459), .E(n18372), .CK(clk), .Q(\RAM<17><5> )
         );
  EDFFX1 \RAM_reg<17><4>  ( .D(n18455), .E(n18373), .CK(clk), .Q(\RAM<17><4> )
         );
  EDFFX1 \RAM_reg<17><3>  ( .D(n18451), .E(n18372), .CK(clk), .Q(\RAM<17><3> )
         );
  EDFFX1 \RAM_reg<17><2>  ( .D(n18447), .E(n18373), .CK(clk), .Q(\RAM<17><2> )
         );
  EDFFX1 \RAM_reg<17><1>  ( .D(n18443), .E(n18372), .CK(clk), .Q(\RAM<17><1> )
         );
  EDFFX1 \RAM_reg<17><0>  ( .D(n18439), .E(n18373), .CK(clk), .Q(\RAM<17><0> )
         );
  EDFFX1 \RAM_reg<9><31>  ( .D(n18564), .E(n18291), .CK(clk), .Q(\RAM<9><31> )
         );
  EDFFX1 \RAM_reg<9><30>  ( .D(n18560), .E(n18291), .CK(clk), .Q(\RAM<9><30> )
         );
  EDFFX1 \RAM_reg<9><29>  ( .D(n18556), .E(n18291), .CK(clk), .Q(\RAM<9><29> )
         );
  EDFFX1 \RAM_reg<9><28>  ( .D(n18552), .E(n18291), .CK(clk), .Q(\RAM<9><28> )
         );
  EDFFX1 \RAM_reg<9><27>  ( .D(n18548), .E(n18291), .CK(clk), .Q(\RAM<9><27> )
         );
  EDFFX1 \RAM_reg<9><26>  ( .D(n18544), .E(n18291), .CK(clk), .Q(\RAM<9><26> )
         );
  EDFFX1 \RAM_reg<9><25>  ( .D(n18540), .E(n18291), .CK(clk), .Q(\RAM<9><25> )
         );
  EDFFX1 \RAM_reg<9><24>  ( .D(n18536), .E(n18291), .CK(clk), .Q(\RAM<9><24> )
         );
  EDFFX1 \RAM_reg<9><23>  ( .D(n18532), .E(n18291), .CK(clk), .Q(\RAM<9><23> )
         );
  EDFFX1 \RAM_reg<9><22>  ( .D(n18528), .E(n18291), .CK(clk), .Q(\RAM<9><22> )
         );
  EDFFX1 \RAM_reg<9><21>  ( .D(n18524), .E(n18291), .CK(clk), .Q(\RAM<9><21> )
         );
  EDFFX1 \RAM_reg<9><20>  ( .D(n18520), .E(n18291), .CK(clk), .Q(\RAM<9><20> )
         );
  EDFFX1 \RAM_reg<9><19>  ( .D(n18516), .E(n18292), .CK(clk), .Q(\RAM<9><19> )
         );
  EDFFX1 \RAM_reg<9><18>  ( .D(n18512), .E(n18292), .CK(clk), .Q(\RAM<9><18> )
         );
  EDFFX1 \RAM_reg<9><17>  ( .D(n18508), .E(n18292), .CK(clk), .Q(\RAM<9><17> )
         );
  EDFFX1 \RAM_reg<9><16>  ( .D(n18504), .E(n18292), .CK(clk), .Q(\RAM<9><16> )
         );
  EDFFX1 \RAM_reg<9><15>  ( .D(n18500), .E(n18292), .CK(clk), .Q(\RAM<9><15> )
         );
  EDFFX1 \RAM_reg<9><14>  ( .D(n18496), .E(n18292), .CK(clk), .Q(\RAM<9><14> )
         );
  EDFFX1 \RAM_reg<9><13>  ( .D(n18492), .E(n18292), .CK(clk), .Q(\RAM<9><13> )
         );
  EDFFX1 \RAM_reg<9><12>  ( .D(n18488), .E(n18292), .CK(clk), .Q(\RAM<9><12> )
         );
  EDFFX1 \RAM_reg<9><11>  ( .D(n18484), .E(n18292), .CK(clk), .Q(\RAM<9><11> )
         );
  EDFFX1 \RAM_reg<9><10>  ( .D(n18480), .E(n18292), .CK(clk), .Q(\RAM<9><10> )
         );
  EDFFX1 \RAM_reg<9><9>  ( .D(n18476), .E(n18292), .CK(clk), .Q(\RAM<9><9> )
         );
  EDFFX1 \RAM_reg<9><8>  ( .D(n18472), .E(n18292), .CK(clk), .Q(\RAM<9><8> )
         );
  EDFFX1 \RAM_reg<9><7>  ( .D(n18468), .E(n3573), .CK(clk), .Q(\RAM<9><7> ) );
  EDFFX1 \RAM_reg<9><6>  ( .D(n18464), .E(n3573), .CK(clk), .Q(\RAM<9><6> ) );
  EDFFX1 \RAM_reg<9><5>  ( .D(n18460), .E(n18291), .CK(clk), .Q(\RAM<9><5> )
         );
  EDFFX1 \RAM_reg<9><4>  ( .D(n18456), .E(n18292), .CK(clk), .Q(\RAM<9><4> )
         );
  EDFFX1 \RAM_reg<9><3>  ( .D(n18452), .E(n18291), .CK(clk), .Q(\RAM<9><3> )
         );
  EDFFX1 \RAM_reg<9><2>  ( .D(n18448), .E(n18292), .CK(clk), .Q(\RAM<9><2> )
         );
  EDFFX1 \RAM_reg<9><1>  ( .D(n18444), .E(n18291), .CK(clk), .Q(\RAM<9><1> )
         );
  EDFFX1 \RAM_reg<9><0>  ( .D(n18440), .E(n18292), .CK(clk), .Q(\RAM<9><0> )
         );
  EDFFX1 \RAM_reg<1><31>  ( .D(n18562), .E(n18297), .CK(clk), .Q(\RAM<1><31> )
         );
  EDFFX1 \RAM_reg<1><30>  ( .D(n18558), .E(n18297), .CK(clk), .Q(\RAM<1><30> )
         );
  EDFFX1 \RAM_reg<1><29>  ( .D(n18554), .E(n18297), .CK(clk), .Q(\RAM<1><29> )
         );
  EDFFX1 \RAM_reg<1><28>  ( .D(n18550), .E(n18297), .CK(clk), .Q(\RAM<1><28> )
         );
  EDFFX1 \RAM_reg<1><27>  ( .D(n18546), .E(n18297), .CK(clk), .Q(\RAM<1><27> )
         );
  EDFFX1 \RAM_reg<1><26>  ( .D(n18542), .E(n18297), .CK(clk), .Q(\RAM<1><26> )
         );
  EDFFX1 \RAM_reg<1><25>  ( .D(n18538), .E(n18297), .CK(clk), .Q(\RAM<1><25> )
         );
  EDFFX1 \RAM_reg<1><24>  ( .D(n18534), .E(n18297), .CK(clk), .Q(\RAM<1><24> )
         );
  EDFFX1 \RAM_reg<1><23>  ( .D(n18530), .E(n18297), .CK(clk), .Q(\RAM<1><23> )
         );
  EDFFX1 \RAM_reg<1><22>  ( .D(n18526), .E(n18297), .CK(clk), .Q(\RAM<1><22> )
         );
  EDFFX1 \RAM_reg<1><21>  ( .D(n18522), .E(n18297), .CK(clk), .Q(\RAM<1><21> )
         );
  EDFFX1 \RAM_reg<1><20>  ( .D(n18518), .E(n18297), .CK(clk), .Q(\RAM<1><20> )
         );
  EDFFX1 \RAM_reg<1><19>  ( .D(n18514), .E(n18298), .CK(clk), .Q(\RAM<1><19> )
         );
  EDFFX1 \RAM_reg<1><18>  ( .D(n18510), .E(n18298), .CK(clk), .Q(\RAM<1><18> )
         );
  EDFFX1 \RAM_reg<1><17>  ( .D(n18506), .E(n18298), .CK(clk), .Q(\RAM<1><17> )
         );
  EDFFX1 \RAM_reg<1><16>  ( .D(n18502), .E(n18298), .CK(clk), .Q(\RAM<1><16> )
         );
  EDFFX1 \RAM_reg<1><15>  ( .D(n18498), .E(n18298), .CK(clk), .Q(\RAM<1><15> )
         );
  EDFFX1 \RAM_reg<1><14>  ( .D(n18494), .E(n18298), .CK(clk), .Q(\RAM<1><14> )
         );
  EDFFX1 \RAM_reg<1><13>  ( .D(n18490), .E(n18298), .CK(clk), .Q(\RAM<1><13> )
         );
  EDFFX1 \RAM_reg<1><12>  ( .D(n18486), .E(n18298), .CK(clk), .Q(\RAM<1><12> )
         );
  EDFFX1 \RAM_reg<1><11>  ( .D(n18482), .E(n18298), .CK(clk), .Q(\RAM<1><11> )
         );
  EDFFX1 \RAM_reg<1><10>  ( .D(n18478), .E(n18298), .CK(clk), .Q(\RAM<1><10> )
         );
  EDFFX1 \RAM_reg<1><9>  ( .D(n18474), .E(n18298), .CK(clk), .Q(\RAM<1><9> )
         );
  EDFFX1 \RAM_reg<1><8>  ( .D(n18470), .E(n18298), .CK(clk), .Q(\RAM<1><8> )
         );
  EDFFX1 \RAM_reg<1><7>  ( .D(n18466), .E(n3571), .CK(clk), .Q(\RAM<1><7> ) );
  EDFFX1 \RAM_reg<1><6>  ( .D(n18462), .E(n3571), .CK(clk), .Q(\RAM<1><6> ) );
  EDFFX1 \RAM_reg<1><5>  ( .D(n18458), .E(n18297), .CK(clk), .Q(\RAM<1><5> )
         );
  EDFFX1 \RAM_reg<1><4>  ( .D(n18454), .E(n18298), .CK(clk), .Q(\RAM<1><4> )
         );
  EDFFX1 \RAM_reg<1><3>  ( .D(n18450), .E(n18297), .CK(clk), .Q(\RAM<1><3> )
         );
  EDFFX1 \RAM_reg<1><2>  ( .D(n18446), .E(n18298), .CK(clk), .Q(\RAM<1><2> )
         );
  EDFFX1 \RAM_reg<1><1>  ( .D(n18442), .E(n18297), .CK(clk), .Q(\RAM<1><1> )
         );
  EDFFX1 \RAM_reg<1><0>  ( .D(n18438), .E(n18298), .CK(clk), .Q(\RAM<1><0> )
         );
  EDFFX1 \RAM_reg<60><31>  ( .D(n18563), .E(n18270), .CK(clk), .Q(
        \RAM<60><31> ) );
  EDFFX1 \RAM_reg<60><30>  ( .D(n18559), .E(n18270), .CK(clk), .Q(
        \RAM<60><30> ) );
  EDFFX1 \RAM_reg<60><29>  ( .D(n18555), .E(n18270), .CK(clk), .Q(
        \RAM<60><29> ) );
  EDFFX1 \RAM_reg<60><28>  ( .D(n18551), .E(n18270), .CK(clk), .Q(
        \RAM<60><28> ) );
  EDFFX1 \RAM_reg<60><27>  ( .D(n18547), .E(n18270), .CK(clk), .Q(
        \RAM<60><27> ) );
  EDFFX1 \RAM_reg<60><26>  ( .D(n18543), .E(n18270), .CK(clk), .Q(
        \RAM<60><26> ) );
  EDFFX1 \RAM_reg<60><25>  ( .D(n18539), .E(n18270), .CK(clk), .Q(
        \RAM<60><25> ) );
  EDFFX1 \RAM_reg<60><24>  ( .D(n18535), .E(n18270), .CK(clk), .Q(
        \RAM<60><24> ) );
  EDFFX1 \RAM_reg<60><23>  ( .D(n18531), .E(n18270), .CK(clk), .Q(
        \RAM<60><23> ) );
  EDFFX1 \RAM_reg<60><22>  ( .D(n18527), .E(n18270), .CK(clk), .Q(
        \RAM<60><22> ) );
  EDFFX1 \RAM_reg<60><21>  ( .D(n18523), .E(n18270), .CK(clk), .Q(
        \RAM<60><21> ) );
  EDFFX1 \RAM_reg<60><20>  ( .D(n18519), .E(n18270), .CK(clk), .Q(
        \RAM<60><20> ) );
  EDFFX1 \RAM_reg<60><19>  ( .D(n18515), .E(n18271), .CK(clk), .Q(
        \RAM<60><19> ) );
  EDFFX1 \RAM_reg<60><18>  ( .D(n18511), .E(n18271), .CK(clk), .Q(
        \RAM<60><18> ) );
  EDFFX1 \RAM_reg<60><17>  ( .D(n18507), .E(n18271), .CK(clk), .Q(
        \RAM<60><17> ) );
  EDFFX1 \RAM_reg<60><16>  ( .D(n18503), .E(n18271), .CK(clk), .Q(
        \RAM<60><16> ) );
  EDFFX1 \RAM_reg<60><15>  ( .D(n18499), .E(n18271), .CK(clk), .Q(
        \RAM<60><15> ) );
  EDFFX1 \RAM_reg<60><14>  ( .D(n18495), .E(n18271), .CK(clk), .Q(
        \RAM<60><14> ) );
  EDFFX1 \RAM_reg<60><13>  ( .D(n18491), .E(n18271), .CK(clk), .Q(
        \RAM<60><13> ) );
  EDFFX1 \RAM_reg<60><12>  ( .D(n18487), .E(n18271), .CK(clk), .Q(
        \RAM<60><12> ) );
  EDFFX1 \RAM_reg<60><11>  ( .D(n18483), .E(n18271), .CK(clk), .Q(
        \RAM<60><11> ) );
  EDFFX1 \RAM_reg<60><10>  ( .D(n18479), .E(n18271), .CK(clk), .Q(
        \RAM<60><10> ) );
  EDFFX1 \RAM_reg<60><9>  ( .D(n18475), .E(n18271), .CK(clk), .Q(\RAM<60><9> )
         );
  EDFFX1 \RAM_reg<60><8>  ( .D(n18471), .E(n18271), .CK(clk), .Q(\RAM<60><8> )
         );
  EDFFX1 \RAM_reg<60><7>  ( .D(n18467), .E(n3581), .CK(clk), .Q(\RAM<60><7> )
         );
  EDFFX1 \RAM_reg<60><6>  ( .D(n18463), .E(n3581), .CK(clk), .Q(\RAM<60><6> )
         );
  EDFFX1 \RAM_reg<60><5>  ( .D(n18459), .E(n18270), .CK(clk), .Q(\RAM<60><5> )
         );
  EDFFX1 \RAM_reg<60><4>  ( .D(n18455), .E(n18271), .CK(clk), .Q(\RAM<60><4> )
         );
  EDFFX1 \RAM_reg<60><3>  ( .D(n18451), .E(n18270), .CK(clk), .Q(\RAM<60><3> )
         );
  EDFFX1 \RAM_reg<60><2>  ( .D(n18447), .E(n18271), .CK(clk), .Q(\RAM<60><2> )
         );
  EDFFX1 \RAM_reg<60><1>  ( .D(n18443), .E(n18270), .CK(clk), .Q(\RAM<60><1> )
         );
  EDFFX1 \RAM_reg<60><0>  ( .D(n18439), .E(n18271), .CK(clk), .Q(\RAM<60><0> )
         );
  EDFFX1 \RAM_reg<56><31>  ( .D(n18564), .E(n18324), .CK(clk), .Q(
        \RAM<56><31> ) );
  EDFFX1 \RAM_reg<56><30>  ( .D(n18560), .E(n18324), .CK(clk), .Q(
        \RAM<56><30> ) );
  EDFFX1 \RAM_reg<56><29>  ( .D(n18556), .E(n18324), .CK(clk), .Q(
        \RAM<56><29> ) );
  EDFFX1 \RAM_reg<56><28>  ( .D(n18552), .E(n18324), .CK(clk), .Q(
        \RAM<56><28> ) );
  EDFFX1 \RAM_reg<56><27>  ( .D(n18548), .E(n18324), .CK(clk), .Q(
        \RAM<56><27> ) );
  EDFFX1 \RAM_reg<56><26>  ( .D(n18544), .E(n18324), .CK(clk), .Q(
        \RAM<56><26> ) );
  EDFFX1 \RAM_reg<56><25>  ( .D(n18540), .E(n18324), .CK(clk), .Q(
        \RAM<56><25> ) );
  EDFFX1 \RAM_reg<56><24>  ( .D(n18536), .E(n18324), .CK(clk), .Q(
        \RAM<56><24> ) );
  EDFFX1 \RAM_reg<56><23>  ( .D(n18532), .E(n18324), .CK(clk), .Q(
        \RAM<56><23> ) );
  EDFFX1 \RAM_reg<56><22>  ( .D(n18528), .E(n18324), .CK(clk), .Q(
        \RAM<56><22> ) );
  EDFFX1 \RAM_reg<56><21>  ( .D(n18524), .E(n18324), .CK(clk), .Q(
        \RAM<56><21> ) );
  EDFFX1 \RAM_reg<56><20>  ( .D(n18520), .E(n18324), .CK(clk), .Q(
        \RAM<56><20> ) );
  EDFFX1 \RAM_reg<56><19>  ( .D(n18516), .E(n18325), .CK(clk), .Q(
        \RAM<56><19> ) );
  EDFFX1 \RAM_reg<56><18>  ( .D(n18512), .E(n18325), .CK(clk), .Q(
        \RAM<56><18> ) );
  EDFFX1 \RAM_reg<56><17>  ( .D(n18508), .E(n18325), .CK(clk), .Q(
        \RAM<56><17> ) );
  EDFFX1 \RAM_reg<56><16>  ( .D(n18504), .E(n18325), .CK(clk), .Q(
        \RAM<56><16> ) );
  EDFFX1 \RAM_reg<56><15>  ( .D(n18500), .E(n18325), .CK(clk), .Q(
        \RAM<56><15> ) );
  EDFFX1 \RAM_reg<56><14>  ( .D(n18496), .E(n18325), .CK(clk), .Q(
        \RAM<56><14> ) );
  EDFFX1 \RAM_reg<56><13>  ( .D(n18492), .E(n18325), .CK(clk), .Q(
        \RAM<56><13> ) );
  EDFFX1 \RAM_reg<56><12>  ( .D(n18488), .E(n18325), .CK(clk), .Q(
        \RAM<56><12> ) );
  EDFFX1 \RAM_reg<56><11>  ( .D(n18484), .E(n18325), .CK(clk), .Q(
        \RAM<56><11> ) );
  EDFFX1 \RAM_reg<56><10>  ( .D(n18480), .E(n18325), .CK(clk), .Q(
        \RAM<56><10> ) );
  EDFFX1 \RAM_reg<56><9>  ( .D(n18476), .E(n18325), .CK(clk), .Q(\RAM<56><9> )
         );
  EDFFX1 \RAM_reg<56><8>  ( .D(n18472), .E(n18325), .CK(clk), .Q(\RAM<56><8> )
         );
  EDFFX1 \RAM_reg<56><7>  ( .D(n18468), .E(n3557), .CK(clk), .Q(\RAM<56><7> )
         );
  EDFFX1 \RAM_reg<56><6>  ( .D(n18464), .E(n3557), .CK(clk), .Q(\RAM<56><6> )
         );
  EDFFX1 \RAM_reg<56><5>  ( .D(n18460), .E(n18324), .CK(clk), .Q(\RAM<56><5> )
         );
  EDFFX1 \RAM_reg<56><4>  ( .D(n18456), .E(n18325), .CK(clk), .Q(\RAM<56><4> )
         );
  EDFFX1 \RAM_reg<56><3>  ( .D(n18452), .E(n18324), .CK(clk), .Q(\RAM<56><3> )
         );
  EDFFX1 \RAM_reg<56><2>  ( .D(n18448), .E(n18325), .CK(clk), .Q(\RAM<56><2> )
         );
  EDFFX1 \RAM_reg<56><1>  ( .D(n18444), .E(n18324), .CK(clk), .Q(\RAM<56><1> )
         );
  EDFFX1 \RAM_reg<56><0>  ( .D(n18440), .E(n18325), .CK(clk), .Q(\RAM<56><0> )
         );
  EDFFX1 \RAM_reg<52><31>  ( .D(n18562), .E(n18342), .CK(clk), .Q(
        \RAM<52><31> ) );
  EDFFX1 \RAM_reg<52><30>  ( .D(n18558), .E(n18342), .CK(clk), .Q(
        \RAM<52><30> ) );
  EDFFX1 \RAM_reg<52><29>  ( .D(n18554), .E(n18342), .CK(clk), .Q(
        \RAM<52><29> ) );
  EDFFX1 \RAM_reg<52><28>  ( .D(n18550), .E(n18342), .CK(clk), .Q(
        \RAM<52><28> ) );
  EDFFX1 \RAM_reg<52><27>  ( .D(n18546), .E(n18342), .CK(clk), .Q(
        \RAM<52><27> ) );
  EDFFX1 \RAM_reg<52><26>  ( .D(n18542), .E(n18342), .CK(clk), .Q(
        \RAM<52><26> ) );
  EDFFX1 \RAM_reg<52><25>  ( .D(n18538), .E(n18342), .CK(clk), .Q(
        \RAM<52><25> ) );
  EDFFX1 \RAM_reg<52><24>  ( .D(n18534), .E(n18342), .CK(clk), .Q(
        \RAM<52><24> ) );
  EDFFX1 \RAM_reg<52><23>  ( .D(n18530), .E(n18342), .CK(clk), .Q(
        \RAM<52><23> ) );
  EDFFX1 \RAM_reg<52><22>  ( .D(n18526), .E(n18342), .CK(clk), .Q(
        \RAM<52><22> ) );
  EDFFX1 \RAM_reg<52><21>  ( .D(n18522), .E(n18342), .CK(clk), .Q(
        \RAM<52><21> ) );
  EDFFX1 \RAM_reg<52><20>  ( .D(n18518), .E(n18342), .CK(clk), .Q(
        \RAM<52><20> ) );
  EDFFX1 \RAM_reg<52><19>  ( .D(n18514), .E(n18343), .CK(clk), .Q(
        \RAM<52><19> ) );
  EDFFX1 \RAM_reg<52><18>  ( .D(n18510), .E(n18343), .CK(clk), .Q(
        \RAM<52><18> ) );
  EDFFX1 \RAM_reg<52><17>  ( .D(n18506), .E(n18343), .CK(clk), .Q(
        \RAM<52><17> ) );
  EDFFX1 \RAM_reg<52><16>  ( .D(n18502), .E(n18343), .CK(clk), .Q(
        \RAM<52><16> ) );
  EDFFX1 \RAM_reg<52><15>  ( .D(n18498), .E(n18343), .CK(clk), .Q(
        \RAM<52><15> ) );
  EDFFX1 \RAM_reg<52><14>  ( .D(n18494), .E(n18343), .CK(clk), .Q(
        \RAM<52><14> ) );
  EDFFX1 \RAM_reg<52><13>  ( .D(n18490), .E(n18343), .CK(clk), .Q(
        \RAM<52><13> ) );
  EDFFX1 \RAM_reg<52><12>  ( .D(n18486), .E(n18343), .CK(clk), .Q(
        \RAM<52><12> ) );
  EDFFX1 \RAM_reg<52><11>  ( .D(n18482), .E(n18343), .CK(clk), .Q(
        \RAM<52><11> ) );
  EDFFX1 \RAM_reg<52><10>  ( .D(n18478), .E(n18343), .CK(clk), .Q(
        \RAM<52><10> ) );
  EDFFX1 \RAM_reg<52><9>  ( .D(n18474), .E(n18343), .CK(clk), .Q(\RAM<52><9> )
         );
  EDFFX1 \RAM_reg<52><8>  ( .D(n18470), .E(n18343), .CK(clk), .Q(\RAM<52><8> )
         );
  EDFFX1 \RAM_reg<52><7>  ( .D(n18466), .E(n3551), .CK(clk), .Q(\RAM<52><7> )
         );
  EDFFX1 \RAM_reg<52><6>  ( .D(n18462), .E(n3551), .CK(clk), .Q(\RAM<52><6> )
         );
  EDFFX1 \RAM_reg<52><5>  ( .D(n18458), .E(n18342), .CK(clk), .Q(\RAM<52><5> )
         );
  EDFFX1 \RAM_reg<52><4>  ( .D(n18454), .E(n18343), .CK(clk), .Q(\RAM<52><4> )
         );
  EDFFX1 \RAM_reg<52><3>  ( .D(n18450), .E(n18342), .CK(clk), .Q(\RAM<52><3> )
         );
  EDFFX1 \RAM_reg<52><2>  ( .D(n18446), .E(n18343), .CK(clk), .Q(\RAM<52><2> )
         );
  EDFFX1 \RAM_reg<52><1>  ( .D(n18442), .E(n18342), .CK(clk), .Q(\RAM<52><1> )
         );
  EDFFX1 \RAM_reg<52><0>  ( .D(n18438), .E(n18343), .CK(clk), .Q(\RAM<52><0> )
         );
  EDFFX1 \RAM_reg<48><31>  ( .D(n18563), .E(n18381), .CK(clk), .Q(
        \RAM<48><31> ) );
  EDFFX1 \RAM_reg<48><30>  ( .D(n18559), .E(n18381), .CK(clk), .Q(
        \RAM<48><30> ) );
  EDFFX1 \RAM_reg<48><29>  ( .D(n18555), .E(n18381), .CK(clk), .Q(
        \RAM<48><29> ) );
  EDFFX1 \RAM_reg<48><28>  ( .D(n18551), .E(n18381), .CK(clk), .Q(
        \RAM<48><28> ) );
  EDFFX1 \RAM_reg<48><27>  ( .D(n18547), .E(n18381), .CK(clk), .Q(
        \RAM<48><27> ) );
  EDFFX1 \RAM_reg<48><26>  ( .D(n18543), .E(n18381), .CK(clk), .Q(
        \RAM<48><26> ) );
  EDFFX1 \RAM_reg<48><25>  ( .D(n18539), .E(n18381), .CK(clk), .Q(
        \RAM<48><25> ) );
  EDFFX1 \RAM_reg<48><24>  ( .D(n18535), .E(n18381), .CK(clk), .Q(
        \RAM<48><24> ) );
  EDFFX1 \RAM_reg<48><23>  ( .D(n18531), .E(n18381), .CK(clk), .Q(
        \RAM<48><23> ) );
  EDFFX1 \RAM_reg<48><22>  ( .D(n18527), .E(n18381), .CK(clk), .Q(
        \RAM<48><22> ) );
  EDFFX1 \RAM_reg<48><21>  ( .D(n18523), .E(n18381), .CK(clk), .Q(
        \RAM<48><21> ) );
  EDFFX1 \RAM_reg<48><20>  ( .D(n18519), .E(n18381), .CK(clk), .Q(
        \RAM<48><20> ) );
  EDFFX1 \RAM_reg<48><19>  ( .D(n18515), .E(n18382), .CK(clk), .Q(
        \RAM<48><19> ) );
  EDFFX1 \RAM_reg<48><18>  ( .D(n18511), .E(n18382), .CK(clk), .Q(
        \RAM<48><18> ) );
  EDFFX1 \RAM_reg<48><17>  ( .D(n18507), .E(n18382), .CK(clk), .Q(
        \RAM<48><17> ) );
  EDFFX1 \RAM_reg<48><16>  ( .D(n18503), .E(n18382), .CK(clk), .Q(
        \RAM<48><16> ) );
  EDFFX1 \RAM_reg<48><15>  ( .D(n18499), .E(n18382), .CK(clk), .Q(
        \RAM<48><15> ) );
  EDFFX1 \RAM_reg<48><14>  ( .D(n18495), .E(n18382), .CK(clk), .Q(
        \RAM<48><14> ) );
  EDFFX1 \RAM_reg<48><13>  ( .D(n18491), .E(n18382), .CK(clk), .Q(
        \RAM<48><13> ) );
  EDFFX1 \RAM_reg<48><12>  ( .D(n18487), .E(n18382), .CK(clk), .Q(
        \RAM<48><12> ) );
  EDFFX1 \RAM_reg<48><11>  ( .D(n18483), .E(n18382), .CK(clk), .Q(
        \RAM<48><11> ) );
  EDFFX1 \RAM_reg<48><10>  ( .D(n18479), .E(n18382), .CK(clk), .Q(
        \RAM<48><10> ) );
  EDFFX1 \RAM_reg<48><9>  ( .D(n18475), .E(n18382), .CK(clk), .Q(\RAM<48><9> )
         );
  EDFFX1 \RAM_reg<48><8>  ( .D(n18471), .E(n18382), .CK(clk), .Q(\RAM<48><8> )
         );
  EDFFX1 \RAM_reg<48><7>  ( .D(n18467), .E(n3536), .CK(clk), .Q(\RAM<48><7> )
         );
  EDFFX1 \RAM_reg<48><6>  ( .D(n18463), .E(n3536), .CK(clk), .Q(\RAM<48><6> )
         );
  EDFFX1 \RAM_reg<48><5>  ( .D(n18459), .E(n18381), .CK(clk), .Q(\RAM<48><5> )
         );
  EDFFX1 \RAM_reg<48><4>  ( .D(n18455), .E(n18382), .CK(clk), .Q(\RAM<48><4> )
         );
  EDFFX1 \RAM_reg<48><3>  ( .D(n18451), .E(n18381), .CK(clk), .Q(\RAM<48><3> )
         );
  EDFFX1 \RAM_reg<48><2>  ( .D(n18447), .E(n18382), .CK(clk), .Q(\RAM<48><2> )
         );
  EDFFX1 \RAM_reg<48><1>  ( .D(n18443), .E(n18381), .CK(clk), .Q(\RAM<48><1> )
         );
  EDFFX1 \RAM_reg<48><0>  ( .D(n18439), .E(n18382), .CK(clk), .Q(\RAM<48><0> )
         );
  EDFFX1 \RAM_reg<44><31>  ( .D(n18564), .E(n18279), .CK(clk), .Q(
        \RAM<44><31> ) );
  EDFFX1 \RAM_reg<44><30>  ( .D(n18560), .E(n18279), .CK(clk), .Q(
        \RAM<44><30> ) );
  EDFFX1 \RAM_reg<44><29>  ( .D(n18556), .E(n18279), .CK(clk), .Q(
        \RAM<44><29> ) );
  EDFFX1 \RAM_reg<44><28>  ( .D(n18552), .E(n18279), .CK(clk), .Q(
        \RAM<44><28> ) );
  EDFFX1 \RAM_reg<44><27>  ( .D(n18548), .E(n18279), .CK(clk), .Q(
        \RAM<44><27> ) );
  EDFFX1 \RAM_reg<44><26>  ( .D(n18544), .E(n18279), .CK(clk), .Q(
        \RAM<44><26> ) );
  EDFFX1 \RAM_reg<44><25>  ( .D(n18540), .E(n18279), .CK(clk), .Q(
        \RAM<44><25> ) );
  EDFFX1 \RAM_reg<44><24>  ( .D(n18536), .E(n18279), .CK(clk), .Q(
        \RAM<44><24> ) );
  EDFFX1 \RAM_reg<44><23>  ( .D(n18532), .E(n18279), .CK(clk), .Q(
        \RAM<44><23> ) );
  EDFFX1 \RAM_reg<44><22>  ( .D(n18528), .E(n18279), .CK(clk), .Q(
        \RAM<44><22> ) );
  EDFFX1 \RAM_reg<44><21>  ( .D(n18524), .E(n18279), .CK(clk), .Q(
        \RAM<44><21> ) );
  EDFFX1 \RAM_reg<44><20>  ( .D(n18520), .E(n18279), .CK(clk), .Q(
        \RAM<44><20> ) );
  EDFFX1 \RAM_reg<44><19>  ( .D(n18516), .E(n18280), .CK(clk), .Q(
        \RAM<44><19> ) );
  EDFFX1 \RAM_reg<44><18>  ( .D(n18512), .E(n18280), .CK(clk), .Q(
        \RAM<44><18> ) );
  EDFFX1 \RAM_reg<44><17>  ( .D(n18508), .E(n18280), .CK(clk), .Q(
        \RAM<44><17> ) );
  EDFFX1 \RAM_reg<44><16>  ( .D(n18504), .E(n18280), .CK(clk), .Q(
        \RAM<44><16> ) );
  EDFFX1 \RAM_reg<44><15>  ( .D(n18500), .E(n18280), .CK(clk), .Q(
        \RAM<44><15> ) );
  EDFFX1 \RAM_reg<44><14>  ( .D(n18496), .E(n18280), .CK(clk), .Q(
        \RAM<44><14> ) );
  EDFFX1 \RAM_reg<44><13>  ( .D(n18492), .E(n18280), .CK(clk), .Q(
        \RAM<44><13> ) );
  EDFFX1 \RAM_reg<44><12>  ( .D(n18488), .E(n18280), .CK(clk), .Q(
        \RAM<44><12> ) );
  EDFFX1 \RAM_reg<44><11>  ( .D(n18484), .E(n18280), .CK(clk), .Q(
        \RAM<44><11> ) );
  EDFFX1 \RAM_reg<44><10>  ( .D(n18480), .E(n18280), .CK(clk), .Q(
        \RAM<44><10> ) );
  EDFFX1 \RAM_reg<44><9>  ( .D(n18476), .E(n18280), .CK(clk), .Q(\RAM<44><9> )
         );
  EDFFX1 \RAM_reg<44><8>  ( .D(n18472), .E(n18280), .CK(clk), .Q(\RAM<44><8> )
         );
  EDFFX1 \RAM_reg<44><7>  ( .D(n18468), .E(n3578), .CK(clk), .Q(\RAM<44><7> )
         );
  EDFFX1 \RAM_reg<44><6>  ( .D(n18464), .E(n3578), .CK(clk), .Q(\RAM<44><6> )
         );
  EDFFX1 \RAM_reg<44><5>  ( .D(n18460), .E(n18279), .CK(clk), .Q(\RAM<44><5> )
         );
  EDFFX1 \RAM_reg<44><4>  ( .D(n18456), .E(n18280), .CK(clk), .Q(\RAM<44><4> )
         );
  EDFFX1 \RAM_reg<44><3>  ( .D(n18452), .E(n18279), .CK(clk), .Q(\RAM<44><3> )
         );
  EDFFX1 \RAM_reg<44><2>  ( .D(n18448), .E(n18280), .CK(clk), .Q(\RAM<44><2> )
         );
  EDFFX1 \RAM_reg<44><1>  ( .D(n18444), .E(n18279), .CK(clk), .Q(\RAM<44><1> )
         );
  EDFFX1 \RAM_reg<44><0>  ( .D(n18440), .E(n18280), .CK(clk), .Q(\RAM<44><0> )
         );
  EDFFX1 \RAM_reg<40><31>  ( .D(n18562), .E(n18396), .CK(clk), .Q(
        \RAM<40><31> ) );
  EDFFX1 \RAM_reg<40><30>  ( .D(n18558), .E(n18396), .CK(clk), .Q(
        \RAM<40><30> ) );
  EDFFX1 \RAM_reg<40><29>  ( .D(n18554), .E(n18396), .CK(clk), .Q(
        \RAM<40><29> ) );
  EDFFX1 \RAM_reg<40><28>  ( .D(n18550), .E(n18396), .CK(clk), .Q(
        \RAM<40><28> ) );
  EDFFX1 \RAM_reg<40><27>  ( .D(n18546), .E(n18396), .CK(clk), .Q(
        \RAM<40><27> ) );
  EDFFX1 \RAM_reg<40><26>  ( .D(n18542), .E(n18396), .CK(clk), .Q(
        \RAM<40><26> ) );
  EDFFX1 \RAM_reg<40><25>  ( .D(n18538), .E(n18396), .CK(clk), .Q(
        \RAM<40><25> ) );
  EDFFX1 \RAM_reg<40><24>  ( .D(n18534), .E(n18396), .CK(clk), .Q(
        \RAM<40><24> ) );
  EDFFX1 \RAM_reg<40><23>  ( .D(n18530), .E(n18396), .CK(clk), .Q(
        \RAM<40><23> ) );
  EDFFX1 \RAM_reg<40><22>  ( .D(n18526), .E(n18396), .CK(clk), .Q(
        \RAM<40><22> ) );
  EDFFX1 \RAM_reg<40><21>  ( .D(n18522), .E(n18396), .CK(clk), .Q(
        \RAM<40><21> ) );
  EDFFX1 \RAM_reg<40><20>  ( .D(n18518), .E(n18396), .CK(clk), .Q(
        \RAM<40><20> ) );
  EDFFX1 \RAM_reg<40><19>  ( .D(n18514), .E(n18397), .CK(clk), .Q(
        \RAM<40><19> ) );
  EDFFX1 \RAM_reg<40><18>  ( .D(n18510), .E(n18397), .CK(clk), .Q(
        \RAM<40><18> ) );
  EDFFX1 \RAM_reg<40><17>  ( .D(n18506), .E(n18397), .CK(clk), .Q(
        \RAM<40><17> ) );
  EDFFX1 \RAM_reg<40><16>  ( .D(n18502), .E(n18397), .CK(clk), .Q(
        \RAM<40><16> ) );
  EDFFX1 \RAM_reg<40><15>  ( .D(n18498), .E(n18397), .CK(clk), .Q(
        \RAM<40><15> ) );
  EDFFX1 \RAM_reg<40><14>  ( .D(n18494), .E(n18397), .CK(clk), .Q(
        \RAM<40><14> ) );
  EDFFX1 \RAM_reg<40><13>  ( .D(n18490), .E(n18397), .CK(clk), .Q(
        \RAM<40><13> ) );
  EDFFX1 \RAM_reg<40><12>  ( .D(n18486), .E(n18397), .CK(clk), .Q(
        \RAM<40><12> ) );
  EDFFX1 \RAM_reg<40><11>  ( .D(n18482), .E(n18397), .CK(clk), .Q(
        \RAM<40><11> ) );
  EDFFX1 \RAM_reg<40><10>  ( .D(n18478), .E(n18397), .CK(clk), .Q(
        \RAM<40><10> ) );
  EDFFX1 \RAM_reg<40><9>  ( .D(n18474), .E(n18397), .CK(clk), .Q(\RAM<40><9> )
         );
  EDFFX1 \RAM_reg<40><8>  ( .D(n18470), .E(n18397), .CK(clk), .Q(\RAM<40><8> )
         );
  EDFFX1 \RAM_reg<40><7>  ( .D(n18466), .E(n3531), .CK(clk), .Q(\RAM<40><7> )
         );
  EDFFX1 \RAM_reg<40><6>  ( .D(n18462), .E(n3531), .CK(clk), .Q(\RAM<40><6> )
         );
  EDFFX1 \RAM_reg<40><5>  ( .D(n18458), .E(n18396), .CK(clk), .Q(\RAM<40><5> )
         );
  EDFFX1 \RAM_reg<40><4>  ( .D(n18454), .E(n18397), .CK(clk), .Q(\RAM<40><4> )
         );
  EDFFX1 \RAM_reg<40><3>  ( .D(n18450), .E(n18396), .CK(clk), .Q(\RAM<40><3> )
         );
  EDFFX1 \RAM_reg<40><2>  ( .D(n18446), .E(n18397), .CK(clk), .Q(\RAM<40><2> )
         );
  EDFFX1 \RAM_reg<40><1>  ( .D(n18442), .E(n18396), .CK(clk), .Q(\RAM<40><1> )
         );
  EDFFX1 \RAM_reg<40><0>  ( .D(n18438), .E(n18397), .CK(clk), .Q(\RAM<40><0> )
         );
  EDFFX1 \RAM_reg<36><31>  ( .D(n18563), .E(n18315), .CK(clk), .Q(
        \RAM<36><31> ) );
  EDFFX1 \RAM_reg<36><30>  ( .D(n18559), .E(n18315), .CK(clk), .Q(
        \RAM<36><30> ) );
  EDFFX1 \RAM_reg<36><29>  ( .D(n18555), .E(n18315), .CK(clk), .Q(
        \RAM<36><29> ) );
  EDFFX1 \RAM_reg<36><28>  ( .D(n18551), .E(n18315), .CK(clk), .Q(
        \RAM<36><28> ) );
  EDFFX1 \RAM_reg<36><27>  ( .D(n18547), .E(n18315), .CK(clk), .Q(
        \RAM<36><27> ) );
  EDFFX1 \RAM_reg<36><26>  ( .D(n18543), .E(n18315), .CK(clk), .Q(
        \RAM<36><26> ) );
  EDFFX1 \RAM_reg<36><25>  ( .D(n18539), .E(n18315), .CK(clk), .Q(
        \RAM<36><25> ) );
  EDFFX1 \RAM_reg<36><24>  ( .D(n18535), .E(n18315), .CK(clk), .Q(
        \RAM<36><24> ) );
  EDFFX1 \RAM_reg<36><23>  ( .D(n18531), .E(n18315), .CK(clk), .Q(
        \RAM<36><23> ) );
  EDFFX1 \RAM_reg<36><22>  ( .D(n18527), .E(n18315), .CK(clk), .Q(
        \RAM<36><22> ) );
  EDFFX1 \RAM_reg<36><21>  ( .D(n18523), .E(n18315), .CK(clk), .Q(
        \RAM<36><21> ) );
  EDFFX1 \RAM_reg<36><20>  ( .D(n18519), .E(n18315), .CK(clk), .Q(
        \RAM<36><20> ) );
  EDFFX1 \RAM_reg<36><19>  ( .D(n18515), .E(n18316), .CK(clk), .Q(
        \RAM<36><19> ) );
  EDFFX1 \RAM_reg<36><18>  ( .D(n18511), .E(n18316), .CK(clk), .Q(
        \RAM<36><18> ) );
  EDFFX1 \RAM_reg<36><17>  ( .D(n18507), .E(n18316), .CK(clk), .Q(
        \RAM<36><17> ) );
  EDFFX1 \RAM_reg<36><16>  ( .D(n18503), .E(n18316), .CK(clk), .Q(
        \RAM<36><16> ) );
  EDFFX1 \RAM_reg<36><15>  ( .D(n18499), .E(n18316), .CK(clk), .Q(
        \RAM<36><15> ) );
  EDFFX1 \RAM_reg<36><14>  ( .D(n18495), .E(n18316), .CK(clk), .Q(
        \RAM<36><14> ) );
  EDFFX1 \RAM_reg<36><13>  ( .D(n18491), .E(n18316), .CK(clk), .Q(
        \RAM<36><13> ) );
  EDFFX1 \RAM_reg<36><12>  ( .D(n18487), .E(n18316), .CK(clk), .Q(
        \RAM<36><12> ) );
  EDFFX1 \RAM_reg<36><11>  ( .D(n18483), .E(n18316), .CK(clk), .Q(
        \RAM<36><11> ) );
  EDFFX1 \RAM_reg<36><10>  ( .D(n18479), .E(n18316), .CK(clk), .Q(
        \RAM<36><10> ) );
  EDFFX1 \RAM_reg<36><9>  ( .D(n18475), .E(n18316), .CK(clk), .Q(\RAM<36><9> )
         );
  EDFFX1 \RAM_reg<36><8>  ( .D(n18471), .E(n18316), .CK(clk), .Q(\RAM<36><8> )
         );
  EDFFX1 \RAM_reg<36><7>  ( .D(n18467), .E(n3562), .CK(clk), .Q(\RAM<36><7> )
         );
  EDFFX1 \RAM_reg<36><6>  ( .D(n18463), .E(n3562), .CK(clk), .Q(\RAM<36><6> )
         );
  EDFFX1 \RAM_reg<36><5>  ( .D(n18459), .E(n18315), .CK(clk), .Q(\RAM<36><5> )
         );
  EDFFX1 \RAM_reg<36><4>  ( .D(n18455), .E(n18316), .CK(clk), .Q(\RAM<36><4> )
         );
  EDFFX1 \RAM_reg<36><3>  ( .D(n18451), .E(n18315), .CK(clk), .Q(\RAM<36><3> )
         );
  EDFFX1 \RAM_reg<36><2>  ( .D(n18447), .E(n18316), .CK(clk), .Q(\RAM<36><2> )
         );
  EDFFX1 \RAM_reg<36><1>  ( .D(n18443), .E(n18315), .CK(clk), .Q(\RAM<36><1> )
         );
  EDFFX1 \RAM_reg<36><0>  ( .D(n18439), .E(n18316), .CK(clk), .Q(\RAM<36><0> )
         );
  EDFFX1 \RAM_reg<32><31>  ( .D(n18564), .E(n18393), .CK(clk), .Q(
        \RAM<32><31> ) );
  EDFFX1 \RAM_reg<32><30>  ( .D(n18560), .E(n18393), .CK(clk), .Q(
        \RAM<32><30> ) );
  EDFFX1 \RAM_reg<32><29>  ( .D(n18556), .E(n18393), .CK(clk), .Q(
        \RAM<32><29> ) );
  EDFFX1 \RAM_reg<32><28>  ( .D(n18552), .E(n18393), .CK(clk), .Q(
        \RAM<32><28> ) );
  EDFFX1 \RAM_reg<32><27>  ( .D(n18548), .E(n18393), .CK(clk), .Q(
        \RAM<32><27> ) );
  EDFFX1 \RAM_reg<32><26>  ( .D(n18544), .E(n18393), .CK(clk), .Q(
        \RAM<32><26> ) );
  EDFFX1 \RAM_reg<32><25>  ( .D(n18540), .E(n18393), .CK(clk), .Q(
        \RAM<32><25> ) );
  EDFFX1 \RAM_reg<32><24>  ( .D(n18536), .E(n18393), .CK(clk), .Q(
        \RAM<32><24> ) );
  EDFFX1 \RAM_reg<32><23>  ( .D(n18532), .E(n18393), .CK(clk), .Q(
        \RAM<32><23> ) );
  EDFFX1 \RAM_reg<32><22>  ( .D(n18528), .E(n18393), .CK(clk), .Q(
        \RAM<32><22> ) );
  EDFFX1 \RAM_reg<32><21>  ( .D(n18524), .E(n18393), .CK(clk), .Q(
        \RAM<32><21> ) );
  EDFFX1 \RAM_reg<32><20>  ( .D(n18520), .E(n18393), .CK(clk), .Q(
        \RAM<32><20> ) );
  EDFFX1 \RAM_reg<32><19>  ( .D(n18516), .E(n18394), .CK(clk), .Q(
        \RAM<32><19> ) );
  EDFFX1 \RAM_reg<32><18>  ( .D(n18512), .E(n18394), .CK(clk), .Q(
        \RAM<32><18> ) );
  EDFFX1 \RAM_reg<32><17>  ( .D(n18508), .E(n18394), .CK(clk), .Q(
        \RAM<32><17> ) );
  EDFFX1 \RAM_reg<32><16>  ( .D(n18504), .E(n18394), .CK(clk), .Q(
        \RAM<32><16> ) );
  EDFFX1 \RAM_reg<32><15>  ( .D(n18500), .E(n18394), .CK(clk), .Q(
        \RAM<32><15> ) );
  EDFFX1 \RAM_reg<32><14>  ( .D(n18496), .E(n18394), .CK(clk), .Q(
        \RAM<32><14> ) );
  EDFFX1 \RAM_reg<32><13>  ( .D(n18492), .E(n18394), .CK(clk), .Q(
        \RAM<32><13> ) );
  EDFFX1 \RAM_reg<32><12>  ( .D(n18488), .E(n18394), .CK(clk), .Q(
        \RAM<32><12> ) );
  EDFFX1 \RAM_reg<32><11>  ( .D(n18484), .E(n18394), .CK(clk), .Q(
        \RAM<32><11> ) );
  EDFFX1 \RAM_reg<32><10>  ( .D(n18480), .E(n18394), .CK(clk), .Q(
        \RAM<32><10> ) );
  EDFFX1 \RAM_reg<32><9>  ( .D(n18476), .E(n18394), .CK(clk), .Q(\RAM<32><9> )
         );
  EDFFX1 \RAM_reg<32><8>  ( .D(n18472), .E(n18394), .CK(clk), .Q(\RAM<32><8> )
         );
  EDFFX1 \RAM_reg<32><7>  ( .D(n18468), .E(n3532), .CK(clk), .Q(\RAM<32><7> )
         );
  EDFFX1 \RAM_reg<32><6>  ( .D(n18464), .E(n3532), .CK(clk), .Q(\RAM<32><6> )
         );
  EDFFX1 \RAM_reg<32><5>  ( .D(n18460), .E(n18393), .CK(clk), .Q(\RAM<32><5> )
         );
  EDFFX1 \RAM_reg<32><4>  ( .D(n18456), .E(n18394), .CK(clk), .Q(\RAM<32><4> )
         );
  EDFFX1 \RAM_reg<32><3>  ( .D(n18452), .E(n18393), .CK(clk), .Q(\RAM<32><3> )
         );
  EDFFX1 \RAM_reg<32><2>  ( .D(n18448), .E(n18394), .CK(clk), .Q(\RAM<32><2> )
         );
  EDFFX1 \RAM_reg<32><1>  ( .D(n18444), .E(n18393), .CK(clk), .Q(\RAM<32><1> )
         );
  EDFFX1 \RAM_reg<32><0>  ( .D(n18440), .E(n18394), .CK(clk), .Q(\RAM<32><0> )
         );
  EDFFX1 \RAM_reg<28><31>  ( .D(n18564), .E(n18366), .CK(clk), .Q(
        \RAM<28><31> ) );
  EDFFX1 \RAM_reg<28><30>  ( .D(n18560), .E(n18366), .CK(clk), .Q(
        \RAM<28><30> ) );
  EDFFX1 \RAM_reg<28><29>  ( .D(n18556), .E(n18366), .CK(clk), .Q(
        \RAM<28><29> ) );
  EDFFX1 \RAM_reg<28><28>  ( .D(n18552), .E(n18366), .CK(clk), .Q(
        \RAM<28><28> ) );
  EDFFX1 \RAM_reg<28><27>  ( .D(n18548), .E(n18366), .CK(clk), .Q(
        \RAM<28><27> ) );
  EDFFX1 \RAM_reg<28><26>  ( .D(n18544), .E(n18366), .CK(clk), .Q(
        \RAM<28><26> ) );
  EDFFX1 \RAM_reg<28><25>  ( .D(n18540), .E(n18366), .CK(clk), .Q(
        \RAM<28><25> ) );
  EDFFX1 \RAM_reg<28><24>  ( .D(n18536), .E(n18366), .CK(clk), .Q(
        \RAM<28><24> ) );
  EDFFX1 \RAM_reg<28><23>  ( .D(n18532), .E(n18366), .CK(clk), .Q(
        \RAM<28><23> ) );
  EDFFX1 \RAM_reg<28><22>  ( .D(n18528), .E(n18366), .CK(clk), .Q(
        \RAM<28><22> ) );
  EDFFX1 \RAM_reg<28><21>  ( .D(n18524), .E(n18366), .CK(clk), .Q(
        \RAM<28><21> ) );
  EDFFX1 \RAM_reg<28><20>  ( .D(n18520), .E(n18366), .CK(clk), .Q(
        \RAM<28><20> ) );
  EDFFX1 \RAM_reg<28><19>  ( .D(n18516), .E(n18367), .CK(clk), .Q(
        \RAM<28><19> ) );
  EDFFX1 \RAM_reg<28><18>  ( .D(n18512), .E(n18367), .CK(clk), .Q(
        \RAM<28><18> ) );
  EDFFX1 \RAM_reg<28><17>  ( .D(n18508), .E(n18367), .CK(clk), .Q(
        \RAM<28><17> ) );
  EDFFX1 \RAM_reg<28><16>  ( .D(n18504), .E(n18367), .CK(clk), .Q(
        \RAM<28><16> ) );
  EDFFX1 \RAM_reg<28><15>  ( .D(n18500), .E(n18367), .CK(clk), .Q(
        \RAM<28><15> ) );
  EDFFX1 \RAM_reg<28><14>  ( .D(n18496), .E(n18367), .CK(clk), .Q(
        \RAM<28><14> ) );
  EDFFX1 \RAM_reg<28><13>  ( .D(n18492), .E(n18367), .CK(clk), .Q(
        \RAM<28><13> ) );
  EDFFX1 \RAM_reg<28><12>  ( .D(n18488), .E(n18367), .CK(clk), .Q(
        \RAM<28><12> ) );
  EDFFX1 \RAM_reg<28><11>  ( .D(n18484), .E(n18367), .CK(clk), .Q(
        \RAM<28><11> ) );
  EDFFX1 \RAM_reg<28><10>  ( .D(n18480), .E(n18367), .CK(clk), .Q(
        \RAM<28><10> ) );
  EDFFX1 \RAM_reg<28><9>  ( .D(n18476), .E(n18367), .CK(clk), .Q(\RAM<28><9> )
         );
  EDFFX1 \RAM_reg<28><8>  ( .D(n18472), .E(n18367), .CK(clk), .Q(\RAM<28><8> )
         );
  EDFFX1 \RAM_reg<28><7>  ( .D(n18468), .E(n3542), .CK(clk), .Q(\RAM<28><7> )
         );
  EDFFX1 \RAM_reg<28><6>  ( .D(n18464), .E(n3542), .CK(clk), .Q(\RAM<28><6> )
         );
  EDFFX1 \RAM_reg<28><5>  ( .D(n18460), .E(n18366), .CK(clk), .Q(\RAM<28><5> )
         );
  EDFFX1 \RAM_reg<28><4>  ( .D(n18456), .E(n18367), .CK(clk), .Q(\RAM<28><4> )
         );
  EDFFX1 \RAM_reg<28><3>  ( .D(n18452), .E(n18366), .CK(clk), .Q(\RAM<28><3> )
         );
  EDFFX1 \RAM_reg<28><2>  ( .D(n18448), .E(n18367), .CK(clk), .Q(\RAM<28><2> )
         );
  EDFFX1 \RAM_reg<28><1>  ( .D(n18444), .E(n18366), .CK(clk), .Q(\RAM<28><1> )
         );
  EDFFX1 \RAM_reg<28><0>  ( .D(n18440), .E(n18367), .CK(clk), .Q(\RAM<28><0> )
         );
  EDFFX1 \RAM_reg<24><31>  ( .D(n18564), .E(n18429), .CK(clk), .Q(
        \RAM<24><31> ) );
  EDFFX1 \RAM_reg<24><30>  ( .D(n18560), .E(n18429), .CK(clk), .Q(
        \RAM<24><30> ) );
  EDFFX1 \RAM_reg<24><29>  ( .D(n18556), .E(n18429), .CK(clk), .Q(
        \RAM<24><29> ) );
  EDFFX1 \RAM_reg<24><28>  ( .D(n18552), .E(n18429), .CK(clk), .Q(
        \RAM<24><28> ) );
  EDFFX1 \RAM_reg<24><27>  ( .D(n18548), .E(n18429), .CK(clk), .Q(
        \RAM<24><27> ) );
  EDFFX1 \RAM_reg<24><26>  ( .D(n18544), .E(n18429), .CK(clk), .Q(
        \RAM<24><26> ) );
  EDFFX1 \RAM_reg<24><25>  ( .D(n18540), .E(n18429), .CK(clk), .Q(
        \RAM<24><25> ) );
  EDFFX1 \RAM_reg<24><24>  ( .D(n18536), .E(n18429), .CK(clk), .Q(
        \RAM<24><24> ) );
  EDFFX1 \RAM_reg<24><23>  ( .D(n18532), .E(n18429), .CK(clk), .Q(
        \RAM<24><23> ) );
  EDFFX1 \RAM_reg<24><22>  ( .D(n18528), .E(n18429), .CK(clk), .Q(
        \RAM<24><22> ) );
  EDFFX1 \RAM_reg<24><21>  ( .D(n18524), .E(n18429), .CK(clk), .Q(
        \RAM<24><21> ) );
  EDFFX1 \RAM_reg<24><20>  ( .D(n18520), .E(n18429), .CK(clk), .Q(
        \RAM<24><20> ) );
  EDFFX1 \RAM_reg<24><19>  ( .D(n18516), .E(n18430), .CK(clk), .Q(
        \RAM<24><19> ) );
  EDFFX1 \RAM_reg<24><18>  ( .D(n18512), .E(n18430), .CK(clk), .Q(
        \RAM<24><18> ) );
  EDFFX1 \RAM_reg<24><17>  ( .D(n18508), .E(n18430), .CK(clk), .Q(
        \RAM<24><17> ) );
  EDFFX1 \RAM_reg<24><16>  ( .D(n18504), .E(n18430), .CK(clk), .Q(
        \RAM<24><16> ) );
  EDFFX1 \RAM_reg<24><15>  ( .D(n18500), .E(n18430), .CK(clk), .Q(
        \RAM<24><15> ) );
  EDFFX1 \RAM_reg<24><14>  ( .D(n18496), .E(n18430), .CK(clk), .Q(
        \RAM<24><14> ) );
  EDFFX1 \RAM_reg<24><13>  ( .D(n18492), .E(n18430), .CK(clk), .Q(
        \RAM<24><13> ) );
  EDFFX1 \RAM_reg<24><12>  ( .D(n18488), .E(n18430), .CK(clk), .Q(
        \RAM<24><12> ) );
  EDFFX1 \RAM_reg<24><11>  ( .D(n18484), .E(n18430), .CK(clk), .Q(
        \RAM<24><11> ) );
  EDFFX1 \RAM_reg<24><10>  ( .D(n18480), .E(n18430), .CK(clk), .Q(
        \RAM<24><10> ) );
  EDFFX1 \RAM_reg<24><9>  ( .D(n18476), .E(n18430), .CK(clk), .Q(\RAM<24><9> )
         );
  EDFFX1 \RAM_reg<24><8>  ( .D(n18472), .E(n18430), .CK(clk), .Q(\RAM<24><8> )
         );
  EDFFX1 \RAM_reg<24><7>  ( .D(n18468), .E(n3520), .CK(clk), .Q(\RAM<24><7> )
         );
  EDFFX1 \RAM_reg<24><6>  ( .D(n18464), .E(n3520), .CK(clk), .Q(\RAM<24><6> )
         );
  EDFFX1 \RAM_reg<24><5>  ( .D(n18460), .E(n18429), .CK(clk), .Q(\RAM<24><5> )
         );
  EDFFX1 \RAM_reg<24><4>  ( .D(n18456), .E(n18430), .CK(clk), .Q(\RAM<24><4> )
         );
  EDFFX1 \RAM_reg<24><3>  ( .D(n18452), .E(n18429), .CK(clk), .Q(\RAM<24><3> )
         );
  EDFFX1 \RAM_reg<24><2>  ( .D(n18448), .E(n18430), .CK(clk), .Q(\RAM<24><2> )
         );
  EDFFX1 \RAM_reg<24><1>  ( .D(n18444), .E(n18429), .CK(clk), .Q(\RAM<24><1> )
         );
  EDFFX1 \RAM_reg<24><0>  ( .D(n18440), .E(n18430), .CK(clk), .Q(\RAM<24><0> )
         );
  EDFFX1 \RAM_reg<20><31>  ( .D(n18564), .E(n18432), .CK(clk), .Q(
        \RAM<20><31> ) );
  EDFFX1 \RAM_reg<20><30>  ( .D(n18560), .E(n18432), .CK(clk), .Q(
        \RAM<20><30> ) );
  EDFFX1 \RAM_reg<20><29>  ( .D(n18556), .E(n18432), .CK(clk), .Q(
        \RAM<20><29> ) );
  EDFFX1 \RAM_reg<20><28>  ( .D(n18552), .E(n18432), .CK(clk), .Q(
        \RAM<20><28> ) );
  EDFFX1 \RAM_reg<20><27>  ( .D(n18548), .E(n18432), .CK(clk), .Q(
        \RAM<20><27> ) );
  EDFFX1 \RAM_reg<20><26>  ( .D(n18544), .E(n18432), .CK(clk), .Q(
        \RAM<20><26> ) );
  EDFFX1 \RAM_reg<20><25>  ( .D(n18540), .E(n18432), .CK(clk), .Q(
        \RAM<20><25> ) );
  EDFFX1 \RAM_reg<20><24>  ( .D(n18536), .E(n18432), .CK(clk), .Q(
        \RAM<20><24> ) );
  EDFFX1 \RAM_reg<20><23>  ( .D(n18532), .E(n18432), .CK(clk), .Q(
        \RAM<20><23> ) );
  EDFFX1 \RAM_reg<20><22>  ( .D(n18528), .E(n18432), .CK(clk), .Q(
        \RAM<20><22> ) );
  EDFFX1 \RAM_reg<20><21>  ( .D(n18524), .E(n18432), .CK(clk), .Q(
        \RAM<20><21> ) );
  EDFFX1 \RAM_reg<20><20>  ( .D(n18520), .E(n18432), .CK(clk), .Q(
        \RAM<20><20> ) );
  EDFFX1 \RAM_reg<20><19>  ( .D(n18516), .E(n18433), .CK(clk), .Q(
        \RAM<20><19> ) );
  EDFFX1 \RAM_reg<20><18>  ( .D(n18512), .E(n18433), .CK(clk), .Q(
        \RAM<20><18> ) );
  EDFFX1 \RAM_reg<20><17>  ( .D(n18508), .E(n18433), .CK(clk), .Q(
        \RAM<20><17> ) );
  EDFFX1 \RAM_reg<20><16>  ( .D(n18504), .E(n18433), .CK(clk), .Q(
        \RAM<20><16> ) );
  EDFFX1 \RAM_reg<20><15>  ( .D(n18500), .E(n18433), .CK(clk), .Q(
        \RAM<20><15> ) );
  EDFFX1 \RAM_reg<20><14>  ( .D(n18496), .E(n18433), .CK(clk), .Q(
        \RAM<20><14> ) );
  EDFFX1 \RAM_reg<20><13>  ( .D(n18492), .E(n18433), .CK(clk), .Q(
        \RAM<20><13> ) );
  EDFFX1 \RAM_reg<20><12>  ( .D(n18488), .E(n18433), .CK(clk), .Q(
        \RAM<20><12> ) );
  EDFFX1 \RAM_reg<20><11>  ( .D(n18484), .E(n18433), .CK(clk), .Q(
        \RAM<20><11> ) );
  EDFFX1 \RAM_reg<20><10>  ( .D(n18480), .E(n18433), .CK(clk), .Q(
        \RAM<20><10> ) );
  EDFFX1 \RAM_reg<20><9>  ( .D(n18476), .E(n18433), .CK(clk), .Q(\RAM<20><9> )
         );
  EDFFX1 \RAM_reg<20><8>  ( .D(n18472), .E(n18433), .CK(clk), .Q(\RAM<20><8> )
         );
  EDFFX1 \RAM_reg<20><7>  ( .D(n18468), .E(n3519), .CK(clk), .Q(\RAM<20><7> )
         );
  EDFFX1 \RAM_reg<20><6>  ( .D(n18464), .E(n3519), .CK(clk), .Q(\RAM<20><6> )
         );
  EDFFX1 \RAM_reg<20><5>  ( .D(n18460), .E(n18432), .CK(clk), .Q(\RAM<20><5> )
         );
  EDFFX1 \RAM_reg<20><4>  ( .D(n18456), .E(n18433), .CK(clk), .Q(\RAM<20><4> )
         );
  EDFFX1 \RAM_reg<20><3>  ( .D(n18452), .E(n18432), .CK(clk), .Q(\RAM<20><3> )
         );
  EDFFX1 \RAM_reg<20><2>  ( .D(n18448), .E(n18433), .CK(clk), .Q(\RAM<20><2> )
         );
  EDFFX1 \RAM_reg<20><1>  ( .D(n18444), .E(n18432), .CK(clk), .Q(\RAM<20><1> )
         );
  EDFFX1 \RAM_reg<20><0>  ( .D(n18440), .E(n18433), .CK(clk), .Q(\RAM<20><0> )
         );
  EDFFX1 \RAM_reg<16><31>  ( .D(n18564), .E(n18309), .CK(clk), .Q(
        \RAM<16><31> ) );
  EDFFX1 \RAM_reg<16><30>  ( .D(n18560), .E(n18309), .CK(clk), .Q(
        \RAM<16><30> ) );
  EDFFX1 \RAM_reg<16><29>  ( .D(n18556), .E(n18309), .CK(clk), .Q(
        \RAM<16><29> ) );
  EDFFX1 \RAM_reg<16><28>  ( .D(n18552), .E(n18309), .CK(clk), .Q(
        \RAM<16><28> ) );
  EDFFX1 \RAM_reg<16><27>  ( .D(n18548), .E(n18309), .CK(clk), .Q(
        \RAM<16><27> ) );
  EDFFX1 \RAM_reg<16><26>  ( .D(n18544), .E(n18309), .CK(clk), .Q(
        \RAM<16><26> ) );
  EDFFX1 \RAM_reg<16><25>  ( .D(n18540), .E(n18309), .CK(clk), .Q(
        \RAM<16><25> ) );
  EDFFX1 \RAM_reg<16><24>  ( .D(n18536), .E(n18309), .CK(clk), .Q(
        \RAM<16><24> ) );
  EDFFX1 \RAM_reg<16><23>  ( .D(n18532), .E(n18309), .CK(clk), .Q(
        \RAM<16><23> ) );
  EDFFX1 \RAM_reg<16><22>  ( .D(n18528), .E(n18309), .CK(clk), .Q(
        \RAM<16><22> ) );
  EDFFX1 \RAM_reg<16><21>  ( .D(n18524), .E(n18309), .CK(clk), .Q(
        \RAM<16><21> ) );
  EDFFX1 \RAM_reg<16><20>  ( .D(n18520), .E(n18309), .CK(clk), .Q(
        \RAM<16><20> ) );
  EDFFX1 \RAM_reg<16><19>  ( .D(n18516), .E(n18310), .CK(clk), .Q(
        \RAM<16><19> ) );
  EDFFX1 \RAM_reg<16><18>  ( .D(n18512), .E(n18310), .CK(clk), .Q(
        \RAM<16><18> ) );
  EDFFX1 \RAM_reg<16><17>  ( .D(n18508), .E(n18310), .CK(clk), .Q(
        \RAM<16><17> ) );
  EDFFX1 \RAM_reg<16><16>  ( .D(n18504), .E(n18310), .CK(clk), .Q(
        \RAM<16><16> ) );
  EDFFX1 \RAM_reg<16><15>  ( .D(n18500), .E(n18310), .CK(clk), .Q(
        \RAM<16><15> ) );
  EDFFX1 \RAM_reg<16><14>  ( .D(n18496), .E(n18310), .CK(clk), .Q(
        \RAM<16><14> ) );
  EDFFX1 \RAM_reg<16><13>  ( .D(n18492), .E(n18310), .CK(clk), .Q(
        \RAM<16><13> ) );
  EDFFX1 \RAM_reg<16><12>  ( .D(n18488), .E(n18310), .CK(clk), .Q(
        \RAM<16><12> ) );
  EDFFX1 \RAM_reg<16><11>  ( .D(n18484), .E(n18310), .CK(clk), .Q(
        \RAM<16><11> ) );
  EDFFX1 \RAM_reg<16><10>  ( .D(n18480), .E(n18310), .CK(clk), .Q(
        \RAM<16><10> ) );
  EDFFX1 \RAM_reg<16><9>  ( .D(n18476), .E(n18310), .CK(clk), .Q(\RAM<16><9> )
         );
  EDFFX1 \RAM_reg<16><8>  ( .D(n18472), .E(n18310), .CK(clk), .Q(\RAM<16><8> )
         );
  EDFFX1 \RAM_reg<16><7>  ( .D(n18468), .E(n3564), .CK(clk), .Q(\RAM<16><7> )
         );
  EDFFX1 \RAM_reg<16><6>  ( .D(n18464), .E(n3564), .CK(clk), .Q(\RAM<16><6> )
         );
  EDFFX1 \RAM_reg<16><5>  ( .D(n18460), .E(n18309), .CK(clk), .Q(\RAM<16><5> )
         );
  EDFFX1 \RAM_reg<16><4>  ( .D(n18456), .E(n18310), .CK(clk), .Q(\RAM<16><4> )
         );
  EDFFX1 \RAM_reg<16><3>  ( .D(n18452), .E(n18309), .CK(clk), .Q(\RAM<16><3> )
         );
  EDFFX1 \RAM_reg<16><2>  ( .D(n18448), .E(n18310), .CK(clk), .Q(\RAM<16><2> )
         );
  EDFFX1 \RAM_reg<16><1>  ( .D(n18444), .E(n18309), .CK(clk), .Q(\RAM<16><1> )
         );
  EDFFX1 \RAM_reg<16><0>  ( .D(n18440), .E(n18310), .CK(clk), .Q(\RAM<16><0> )
         );
  EDFFX1 \RAM_reg<12><31>  ( .D(n18564), .E(n18273), .CK(clk), .Q(
        \RAM<12><31> ) );
  EDFFX1 \RAM_reg<12><30>  ( .D(n18560), .E(n18273), .CK(clk), .Q(
        \RAM<12><30> ) );
  EDFFX1 \RAM_reg<12><29>  ( .D(n18556), .E(n18273), .CK(clk), .Q(
        \RAM<12><29> ) );
  EDFFX1 \RAM_reg<12><28>  ( .D(n18552), .E(n18273), .CK(clk), .Q(
        \RAM<12><28> ) );
  EDFFX1 \RAM_reg<12><27>  ( .D(n18548), .E(n18273), .CK(clk), .Q(
        \RAM<12><27> ) );
  EDFFX1 \RAM_reg<12><26>  ( .D(n18544), .E(n18273), .CK(clk), .Q(
        \RAM<12><26> ) );
  EDFFX1 \RAM_reg<12><25>  ( .D(n18540), .E(n18273), .CK(clk), .Q(
        \RAM<12><25> ) );
  EDFFX1 \RAM_reg<12><24>  ( .D(n18536), .E(n18273), .CK(clk), .Q(
        \RAM<12><24> ) );
  EDFFX1 \RAM_reg<12><23>  ( .D(n18532), .E(n18273), .CK(clk), .Q(
        \RAM<12><23> ) );
  EDFFX1 \RAM_reg<12><22>  ( .D(n18528), .E(n18273), .CK(clk), .Q(
        \RAM<12><22> ) );
  EDFFX1 \RAM_reg<12><21>  ( .D(n18524), .E(n18273), .CK(clk), .Q(
        \RAM<12><21> ) );
  EDFFX1 \RAM_reg<12><20>  ( .D(n18520), .E(n18273), .CK(clk), .Q(
        \RAM<12><20> ) );
  EDFFX1 \RAM_reg<12><19>  ( .D(n18516), .E(n18274), .CK(clk), .Q(
        \RAM<12><19> ) );
  EDFFX1 \RAM_reg<12><18>  ( .D(n18512), .E(n18274), .CK(clk), .Q(
        \RAM<12><18> ) );
  EDFFX1 \RAM_reg<12><17>  ( .D(n18508), .E(n18274), .CK(clk), .Q(
        \RAM<12><17> ) );
  EDFFX1 \RAM_reg<12><16>  ( .D(n18504), .E(n18274), .CK(clk), .Q(
        \RAM<12><16> ) );
  EDFFX1 \RAM_reg<12><15>  ( .D(n18500), .E(n18274), .CK(clk), .Q(
        \RAM<12><15> ) );
  EDFFX1 \RAM_reg<12><14>  ( .D(n18496), .E(n18274), .CK(clk), .Q(
        \RAM<12><14> ) );
  EDFFX1 \RAM_reg<12><13>  ( .D(n18492), .E(n18274), .CK(clk), .Q(
        \RAM<12><13> ) );
  EDFFX1 \RAM_reg<12><12>  ( .D(n18488), .E(n18274), .CK(clk), .Q(
        \RAM<12><12> ) );
  EDFFX1 \RAM_reg<12><11>  ( .D(n18484), .E(n18274), .CK(clk), .Q(
        \RAM<12><11> ) );
  EDFFX1 \RAM_reg<12><10>  ( .D(n18480), .E(n18274), .CK(clk), .Q(
        \RAM<12><10> ) );
  EDFFX1 \RAM_reg<12><9>  ( .D(n18476), .E(n18274), .CK(clk), .Q(\RAM<12><9> )
         );
  EDFFX1 \RAM_reg<12><8>  ( .D(n18472), .E(n18274), .CK(clk), .Q(\RAM<12><8> )
         );
  EDFFX1 \RAM_reg<12><7>  ( .D(n18468), .E(n3580), .CK(clk), .Q(\RAM<12><7> )
         );
  EDFFX1 \RAM_reg<12><6>  ( .D(n18464), .E(n3580), .CK(clk), .Q(\RAM<12><6> )
         );
  EDFFX1 \RAM_reg<12><5>  ( .D(n18460), .E(n18273), .CK(clk), .Q(\RAM<12><5> )
         );
  EDFFX1 \RAM_reg<12><4>  ( .D(n18456), .E(n18274), .CK(clk), .Q(\RAM<12><4> )
         );
  EDFFX1 \RAM_reg<12><3>  ( .D(n18452), .E(n18273), .CK(clk), .Q(\RAM<12><3> )
         );
  EDFFX1 \RAM_reg<12><2>  ( .D(n18448), .E(n18274), .CK(clk), .Q(\RAM<12><2> )
         );
  EDFFX1 \RAM_reg<12><1>  ( .D(n18444), .E(n18273), .CK(clk), .Q(\RAM<12><1> )
         );
  EDFFX1 \RAM_reg<12><0>  ( .D(n18440), .E(n18274), .CK(clk), .Q(\RAM<12><0> )
         );
  EDFFX1 \RAM_reg<8><31>  ( .D(n18564), .E(n18306), .CK(clk), .Q(\RAM<8><31> )
         );
  EDFFX1 \RAM_reg<8><30>  ( .D(n18560), .E(n18306), .CK(clk), .Q(\RAM<8><30> )
         );
  EDFFX1 \RAM_reg<8><29>  ( .D(n18556), .E(n18306), .CK(clk), .Q(\RAM<8><29> )
         );
  EDFFX1 \RAM_reg<8><28>  ( .D(n18552), .E(n18306), .CK(clk), .Q(\RAM<8><28> )
         );
  EDFFX1 \RAM_reg<8><27>  ( .D(n18548), .E(n18306), .CK(clk), .Q(\RAM<8><27> )
         );
  EDFFX1 \RAM_reg<8><26>  ( .D(n18544), .E(n18306), .CK(clk), .Q(\RAM<8><26> )
         );
  EDFFX1 \RAM_reg<8><25>  ( .D(n18540), .E(n18306), .CK(clk), .Q(\RAM<8><25> )
         );
  EDFFX1 \RAM_reg<8><24>  ( .D(n18536), .E(n18306), .CK(clk), .Q(\RAM<8><24> )
         );
  EDFFX1 \RAM_reg<8><23>  ( .D(n18532), .E(n18306), .CK(clk), .Q(\RAM<8><23> )
         );
  EDFFX1 \RAM_reg<8><22>  ( .D(n18528), .E(n18306), .CK(clk), .Q(\RAM<8><22> )
         );
  EDFFX1 \RAM_reg<8><21>  ( .D(n18524), .E(n18306), .CK(clk), .Q(\RAM<8><21> )
         );
  EDFFX1 \RAM_reg<8><20>  ( .D(n18520), .E(n18306), .CK(clk), .Q(\RAM<8><20> )
         );
  EDFFX1 \RAM_reg<8><19>  ( .D(n18516), .E(n18307), .CK(clk), .Q(\RAM<8><19> )
         );
  EDFFX1 \RAM_reg<8><18>  ( .D(n18512), .E(n18307), .CK(clk), .Q(\RAM<8><18> )
         );
  EDFFX1 \RAM_reg<8><17>  ( .D(n18508), .E(n18307), .CK(clk), .Q(\RAM<8><17> )
         );
  EDFFX1 \RAM_reg<8><16>  ( .D(n18504), .E(n18307), .CK(clk), .Q(\RAM<8><16> )
         );
  EDFFX1 \RAM_reg<8><15>  ( .D(n18500), .E(n18307), .CK(clk), .Q(\RAM<8><15> )
         );
  EDFFX1 \RAM_reg<8><14>  ( .D(n18496), .E(n18307), .CK(clk), .Q(\RAM<8><14> )
         );
  EDFFX1 \RAM_reg<8><13>  ( .D(n18492), .E(n18307), .CK(clk), .Q(\RAM<8><13> )
         );
  EDFFX1 \RAM_reg<8><12>  ( .D(n18488), .E(n18307), .CK(clk), .Q(\RAM<8><12> )
         );
  EDFFX1 \RAM_reg<8><11>  ( .D(n18484), .E(n18307), .CK(clk), .Q(\RAM<8><11> )
         );
  EDFFX1 \RAM_reg<8><10>  ( .D(n18480), .E(n18307), .CK(clk), .Q(\RAM<8><10> )
         );
  EDFFX1 \RAM_reg<8><9>  ( .D(n18476), .E(n18307), .CK(clk), .Q(\RAM<8><9> )
         );
  EDFFX1 \RAM_reg<8><8>  ( .D(n18472), .E(n18307), .CK(clk), .Q(\RAM<8><8> )
         );
  EDFFX1 \RAM_reg<8><7>  ( .D(n18468), .E(n3567), .CK(clk), .Q(\RAM<8><7> ) );
  EDFFX1 \RAM_reg<8><6>  ( .D(n18464), .E(n3567), .CK(clk), .Q(\RAM<8><6> ) );
  EDFFX1 \RAM_reg<8><5>  ( .D(n18460), .E(n18306), .CK(clk), .Q(\RAM<8><5> )
         );
  EDFFX1 \RAM_reg<8><4>  ( .D(n18456), .E(n18307), .CK(clk), .Q(\RAM<8><4> )
         );
  EDFFX1 \RAM_reg<8><3>  ( .D(n18452), .E(n18306), .CK(clk), .Q(\RAM<8><3> )
         );
  EDFFX1 \RAM_reg<8><2>  ( .D(n18448), .E(n18307), .CK(clk), .Q(\RAM<8><2> )
         );
  EDFFX1 \RAM_reg<8><1>  ( .D(n18444), .E(n18306), .CK(clk), .Q(\RAM<8><1> )
         );
  EDFFX1 \RAM_reg<8><0>  ( .D(n18440), .E(n18307), .CK(clk), .Q(\RAM<8><0> )
         );
  EDFFX1 \RAM_reg<4><31>  ( .D(n18564), .E(n18276), .CK(clk), .Q(\RAM<4><31> )
         );
  EDFFX1 \RAM_reg<4><30>  ( .D(n18560), .E(n18276), .CK(clk), .Q(\RAM<4><30> )
         );
  EDFFX1 \RAM_reg<4><29>  ( .D(n18556), .E(n18276), .CK(clk), .Q(\RAM<4><29> )
         );
  EDFFX1 \RAM_reg<4><28>  ( .D(n18552), .E(n18276), .CK(clk), .Q(\RAM<4><28> )
         );
  EDFFX1 \RAM_reg<4><27>  ( .D(n18548), .E(n18276), .CK(clk), .Q(\RAM<4><27> )
         );
  EDFFX1 \RAM_reg<4><26>  ( .D(n18544), .E(n18276), .CK(clk), .Q(\RAM<4><26> )
         );
  EDFFX1 \RAM_reg<4><25>  ( .D(n18540), .E(n18276), .CK(clk), .Q(\RAM<4><25> )
         );
  EDFFX1 \RAM_reg<4><24>  ( .D(n18536), .E(n18276), .CK(clk), .Q(\RAM<4><24> )
         );
  EDFFX1 \RAM_reg<4><23>  ( .D(n18532), .E(n18276), .CK(clk), .Q(\RAM<4><23> )
         );
  EDFFX1 \RAM_reg<4><22>  ( .D(n18528), .E(n18276), .CK(clk), .Q(\RAM<4><22> )
         );
  EDFFX1 \RAM_reg<4><21>  ( .D(n18524), .E(n18276), .CK(clk), .Q(\RAM<4><21> )
         );
  EDFFX1 \RAM_reg<4><20>  ( .D(n18520), .E(n18276), .CK(clk), .Q(\RAM<4><20> )
         );
  EDFFX1 \RAM_reg<4><19>  ( .D(n18516), .E(n18277), .CK(clk), .Q(\RAM<4><19> )
         );
  EDFFX1 \RAM_reg<4><18>  ( .D(n18512), .E(n18277), .CK(clk), .Q(\RAM<4><18> )
         );
  EDFFX1 \RAM_reg<4><17>  ( .D(n18508), .E(n18277), .CK(clk), .Q(\RAM<4><17> )
         );
  EDFFX1 \RAM_reg<4><16>  ( .D(n18504), .E(n18277), .CK(clk), .Q(\RAM<4><16> )
         );
  EDFFX1 \RAM_reg<4><15>  ( .D(n18500), .E(n18277), .CK(clk), .Q(\RAM<4><15> )
         );
  EDFFX1 \RAM_reg<4><14>  ( .D(n18496), .E(n18277), .CK(clk), .Q(\RAM<4><14> )
         );
  EDFFX1 \RAM_reg<4><13>  ( .D(n18492), .E(n18277), .CK(clk), .Q(\RAM<4><13> )
         );
  EDFFX1 \RAM_reg<4><12>  ( .D(n18488), .E(n18277), .CK(clk), .Q(\RAM<4><12> )
         );
  EDFFX1 \RAM_reg<4><11>  ( .D(n18484), .E(n18277), .CK(clk), .Q(\RAM<4><11> )
         );
  EDFFX1 \RAM_reg<4><10>  ( .D(n18480), .E(n18277), .CK(clk), .Q(\RAM<4><10> )
         );
  EDFFX1 \RAM_reg<4><9>  ( .D(n18476), .E(n18277), .CK(clk), .Q(\RAM<4><9> )
         );
  EDFFX1 \RAM_reg<4><8>  ( .D(n18472), .E(n18277), .CK(clk), .Q(\RAM<4><8> )
         );
  EDFFX1 \RAM_reg<4><7>  ( .D(n18468), .E(n3579), .CK(clk), .Q(\RAM<4><7> ) );
  EDFFX1 \RAM_reg<4><6>  ( .D(n18464), .E(n3579), .CK(clk), .Q(\RAM<4><6> ) );
  EDFFX1 \RAM_reg<4><5>  ( .D(n18460), .E(n18276), .CK(clk), .Q(\RAM<4><5> )
         );
  EDFFX1 \RAM_reg<4><4>  ( .D(n18456), .E(n18277), .CK(clk), .Q(\RAM<4><4> )
         );
  EDFFX1 \RAM_reg<4><3>  ( .D(n18452), .E(n18276), .CK(clk), .Q(\RAM<4><3> )
         );
  EDFFX1 \RAM_reg<4><2>  ( .D(n18448), .E(n18277), .CK(clk), .Q(\RAM<4><2> )
         );
  EDFFX1 \RAM_reg<4><1>  ( .D(n18444), .E(n18276), .CK(clk), .Q(\RAM<4><1> )
         );
  EDFFX1 \RAM_reg<4><0>  ( .D(n18440), .E(n18277), .CK(clk), .Q(\RAM<4><0> )
         );
  EDFFX1 \RAM_reg<0><31>  ( .D(n18564), .E(n18333), .CK(clk), .Q(\RAM<0><31> )
         );
  EDFFX1 \RAM_reg<0><30>  ( .D(n18560), .E(n18333), .CK(clk), .Q(\RAM<0><30> )
         );
  EDFFX1 \RAM_reg<0><29>  ( .D(n18556), .E(n18333), .CK(clk), .Q(\RAM<0><29> )
         );
  EDFFX1 \RAM_reg<0><28>  ( .D(n18552), .E(n18333), .CK(clk), .Q(\RAM<0><28> )
         );
  EDFFX1 \RAM_reg<0><27>  ( .D(n18548), .E(n18333), .CK(clk), .Q(\RAM<0><27> )
         );
  EDFFX1 \RAM_reg<0><26>  ( .D(n18544), .E(n18333), .CK(clk), .Q(\RAM<0><26> )
         );
  EDFFX1 \RAM_reg<0><25>  ( .D(n18540), .E(n18333), .CK(clk), .Q(\RAM<0><25> )
         );
  EDFFX1 \RAM_reg<0><24>  ( .D(n18536), .E(n18333), .CK(clk), .Q(\RAM<0><24> )
         );
  EDFFX1 \RAM_reg<0><23>  ( .D(n18532), .E(n18333), .CK(clk), .Q(\RAM<0><23> )
         );
  EDFFX1 \RAM_reg<0><22>  ( .D(n18528), .E(n18333), .CK(clk), .Q(\RAM<0><22> )
         );
  EDFFX1 \RAM_reg<0><21>  ( .D(n18524), .E(n18333), .CK(clk), .Q(\RAM<0><21> )
         );
  EDFFX1 \RAM_reg<0><20>  ( .D(n18520), .E(n18333), .CK(clk), .Q(\RAM<0><20> )
         );
  EDFFX1 \RAM_reg<0><19>  ( .D(n18516), .E(n18334), .CK(clk), .Q(\RAM<0><19> )
         );
  EDFFX1 \RAM_reg<0><18>  ( .D(n18512), .E(n18334), .CK(clk), .Q(\RAM<0><18> )
         );
  EDFFX1 \RAM_reg<0><17>  ( .D(n18508), .E(n18334), .CK(clk), .Q(\RAM<0><17> )
         );
  EDFFX1 \RAM_reg<0><16>  ( .D(n18504), .E(n18334), .CK(clk), .Q(\RAM<0><16> )
         );
  EDFFX1 \RAM_reg<0><15>  ( .D(n18500), .E(n18334), .CK(clk), .Q(\RAM<0><15> )
         );
  EDFFX1 \RAM_reg<0><14>  ( .D(n18496), .E(n18334), .CK(clk), .Q(\RAM<0><14> )
         );
  EDFFX1 \RAM_reg<0><13>  ( .D(n18492), .E(n18334), .CK(clk), .Q(\RAM<0><13> )
         );
  EDFFX1 \RAM_reg<0><12>  ( .D(n18488), .E(n18334), .CK(clk), .Q(\RAM<0><12> )
         );
  EDFFX1 \RAM_reg<0><11>  ( .D(n18484), .E(n18334), .CK(clk), .Q(\RAM<0><11> )
         );
  EDFFX1 \RAM_reg<0><10>  ( .D(n18480), .E(n18334), .CK(clk), .Q(\RAM<0><10> )
         );
  EDFFX1 \RAM_reg<0><9>  ( .D(n18476), .E(n18334), .CK(clk), .Q(\RAM<0><9> )
         );
  EDFFX1 \RAM_reg<0><8>  ( .D(n18472), .E(n18334), .CK(clk), .Q(\RAM<0><8> )
         );
  EDFFX1 \RAM_reg<0><7>  ( .D(n18468), .E(n3554), .CK(clk), .Q(\RAM<0><7> ) );
  EDFFX1 \RAM_reg<0><6>  ( .D(n18464), .E(n3554), .CK(clk), .Q(\RAM<0><6> ) );
  EDFFX1 \RAM_reg<0><5>  ( .D(n18460), .E(n18333), .CK(clk), .Q(\RAM<0><5> )
         );
  EDFFX1 \RAM_reg<0><4>  ( .D(n18456), .E(n18334), .CK(clk), .Q(\RAM<0><4> )
         );
  EDFFX1 \RAM_reg<0><3>  ( .D(n18452), .E(n18333), .CK(clk), .Q(\RAM<0><3> )
         );
  EDFFX1 \RAM_reg<0><2>  ( .D(n18448), .E(n18334), .CK(clk), .Q(\RAM<0><2> )
         );
  EDFFX1 \RAM_reg<0><1>  ( .D(n18444), .E(n18333), .CK(clk), .Q(\RAM<0><1> )
         );
  EDFFX1 \RAM_reg<0><0>  ( .D(n18440), .E(n18334), .CK(clk), .Q(\RAM<0><0> )
         );
  EDFFX1 \RAM_reg<62><31>  ( .D(n18564), .E(n18357), .CK(clk), .Q(
        \RAM<62><31> ) );
  EDFFX1 \RAM_reg<62><30>  ( .D(n18560), .E(n18357), .CK(clk), .Q(
        \RAM<62><30> ) );
  EDFFX1 \RAM_reg<62><29>  ( .D(n18556), .E(n18357), .CK(clk), .Q(
        \RAM<62><29> ) );
  EDFFX1 \RAM_reg<62><28>  ( .D(n18552), .E(n18357), .CK(clk), .Q(
        \RAM<62><28> ) );
  EDFFX1 \RAM_reg<62><27>  ( .D(n18548), .E(n18357), .CK(clk), .Q(
        \RAM<62><27> ) );
  EDFFX1 \RAM_reg<62><26>  ( .D(n18544), .E(n18357), .CK(clk), .Q(
        \RAM<62><26> ) );
  EDFFX1 \RAM_reg<62><25>  ( .D(n18540), .E(n18357), .CK(clk), .Q(
        \RAM<62><25> ) );
  EDFFX1 \RAM_reg<62><24>  ( .D(n18536), .E(n18357), .CK(clk), .Q(
        \RAM<62><24> ) );
  EDFFX1 \RAM_reg<62><23>  ( .D(n18532), .E(n18357), .CK(clk), .Q(
        \RAM<62><23> ) );
  EDFFX1 \RAM_reg<62><22>  ( .D(n18528), .E(n18357), .CK(clk), .Q(
        \RAM<62><22> ) );
  EDFFX1 \RAM_reg<62><21>  ( .D(n18524), .E(n18357), .CK(clk), .Q(
        \RAM<62><21> ) );
  EDFFX1 \RAM_reg<62><20>  ( .D(n18520), .E(n18357), .CK(clk), .Q(
        \RAM<62><20> ) );
  EDFFX1 \RAM_reg<62><19>  ( .D(n18516), .E(n18358), .CK(clk), .Q(
        \RAM<62><19> ) );
  EDFFX1 \RAM_reg<62><18>  ( .D(n18512), .E(n18358), .CK(clk), .Q(
        \RAM<62><18> ) );
  EDFFX1 \RAM_reg<62><17>  ( .D(n18508), .E(n18358), .CK(clk), .Q(
        \RAM<62><17> ) );
  EDFFX1 \RAM_reg<62><16>  ( .D(n18504), .E(n18358), .CK(clk), .Q(
        \RAM<62><16> ) );
  EDFFX1 \RAM_reg<62><15>  ( .D(n18500), .E(n18358), .CK(clk), .Q(
        \RAM<62><15> ) );
  EDFFX1 \RAM_reg<62><14>  ( .D(n18496), .E(n18358), .CK(clk), .Q(
        \RAM<62><14> ) );
  EDFFX1 \RAM_reg<62><13>  ( .D(n18492), .E(n18358), .CK(clk), .Q(
        \RAM<62><13> ) );
  EDFFX1 \RAM_reg<62><12>  ( .D(n18488), .E(n18358), .CK(clk), .Q(
        \RAM<62><12> ) );
  EDFFX1 \RAM_reg<62><11>  ( .D(n18484), .E(n18358), .CK(clk), .Q(
        \RAM<62><11> ) );
  EDFFX1 \RAM_reg<62><10>  ( .D(n18480), .E(n18358), .CK(clk), .Q(
        \RAM<62><10> ) );
  EDFFX1 \RAM_reg<62><9>  ( .D(n18476), .E(n18358), .CK(clk), .Q(\RAM<62><9> )
         );
  EDFFX1 \RAM_reg<62><8>  ( .D(n18472), .E(n18358), .CK(clk), .Q(\RAM<62><8> )
         );
  EDFFX1 \RAM_reg<62><7>  ( .D(n18468), .E(n3545), .CK(clk), .Q(\RAM<62><7> )
         );
  EDFFX1 \RAM_reg<62><6>  ( .D(n18464), .E(n3545), .CK(clk), .Q(\RAM<62><6> )
         );
  EDFFX1 \RAM_reg<62><5>  ( .D(n18460), .E(n18357), .CK(clk), .Q(\RAM<62><5> )
         );
  EDFFX1 \RAM_reg<62><4>  ( .D(n18456), .E(n18358), .CK(clk), .Q(\RAM<62><4> )
         );
  EDFFX1 \RAM_reg<62><3>  ( .D(n18452), .E(n18357), .CK(clk), .Q(\RAM<62><3> )
         );
  EDFFX1 \RAM_reg<62><2>  ( .D(n18448), .E(n18358), .CK(clk), .Q(\RAM<62><2> )
         );
  EDFFX1 \RAM_reg<62><1>  ( .D(n18444), .E(n18357), .CK(clk), .Q(\RAM<62><1> )
         );
  EDFFX1 \RAM_reg<62><0>  ( .D(n18440), .E(n18358), .CK(clk), .Q(\RAM<62><0> )
         );
  EDFFX1 \RAM_reg<54><31>  ( .D(n18564), .E(n18348), .CK(clk), .Q(
        \RAM<54><31> ) );
  EDFFX1 \RAM_reg<54><30>  ( .D(n18560), .E(n18348), .CK(clk), .Q(
        \RAM<54><30> ) );
  EDFFX1 \RAM_reg<54><29>  ( .D(n18556), .E(n18348), .CK(clk), .Q(
        \RAM<54><29> ) );
  EDFFX1 \RAM_reg<54><28>  ( .D(n18552), .E(n18348), .CK(clk), .Q(
        \RAM<54><28> ) );
  EDFFX1 \RAM_reg<54><27>  ( .D(n18548), .E(n18348), .CK(clk), .Q(
        \RAM<54><27> ) );
  EDFFX1 \RAM_reg<54><26>  ( .D(n18544), .E(n18348), .CK(clk), .Q(
        \RAM<54><26> ) );
  EDFFX1 \RAM_reg<54><25>  ( .D(n18540), .E(n18348), .CK(clk), .Q(
        \RAM<54><25> ) );
  EDFFX1 \RAM_reg<54><24>  ( .D(n18536), .E(n18348), .CK(clk), .Q(
        \RAM<54><24> ) );
  EDFFX1 \RAM_reg<54><23>  ( .D(n18532), .E(n18348), .CK(clk), .Q(
        \RAM<54><23> ) );
  EDFFX1 \RAM_reg<54><22>  ( .D(n18528), .E(n18348), .CK(clk), .Q(
        \RAM<54><22> ) );
  EDFFX1 \RAM_reg<54><21>  ( .D(n18524), .E(n18348), .CK(clk), .Q(
        \RAM<54><21> ) );
  EDFFX1 \RAM_reg<54><20>  ( .D(n18520), .E(n18348), .CK(clk), .Q(
        \RAM<54><20> ) );
  EDFFX1 \RAM_reg<54><19>  ( .D(n18516), .E(n18349), .CK(clk), .Q(
        \RAM<54><19> ) );
  EDFFX1 \RAM_reg<54><18>  ( .D(n18512), .E(n18349), .CK(clk), .Q(
        \RAM<54><18> ) );
  EDFFX1 \RAM_reg<54><17>  ( .D(n18508), .E(n18349), .CK(clk), .Q(
        \RAM<54><17> ) );
  EDFFX1 \RAM_reg<54><16>  ( .D(n18504), .E(n18349), .CK(clk), .Q(
        \RAM<54><16> ) );
  EDFFX1 \RAM_reg<54><15>  ( .D(n18500), .E(n18349), .CK(clk), .Q(
        \RAM<54><15> ) );
  EDFFX1 \RAM_reg<54><14>  ( .D(n18496), .E(n18349), .CK(clk), .Q(
        \RAM<54><14> ) );
  EDFFX1 \RAM_reg<54><13>  ( .D(n18492), .E(n18349), .CK(clk), .Q(
        \RAM<54><13> ) );
  EDFFX1 \RAM_reg<54><12>  ( .D(n18488), .E(n18349), .CK(clk), .Q(
        \RAM<54><12> ) );
  EDFFX1 \RAM_reg<54><11>  ( .D(n18484), .E(n18349), .CK(clk), .Q(
        \RAM<54><11> ) );
  EDFFX1 \RAM_reg<54><10>  ( .D(n18480), .E(n18349), .CK(clk), .Q(
        \RAM<54><10> ) );
  EDFFX1 \RAM_reg<54><9>  ( .D(n18476), .E(n18349), .CK(clk), .Q(\RAM<54><9> )
         );
  EDFFX1 \RAM_reg<54><8>  ( .D(n18472), .E(n18349), .CK(clk), .Q(\RAM<54><8> )
         );
  EDFFX1 \RAM_reg<54><7>  ( .D(n18468), .E(n3549), .CK(clk), .Q(\RAM<54><7> )
         );
  EDFFX1 \RAM_reg<54><6>  ( .D(n18464), .E(n3549), .CK(clk), .Q(\RAM<54><6> )
         );
  EDFFX1 \RAM_reg<54><5>  ( .D(n18460), .E(n18348), .CK(clk), .Q(\RAM<54><5> )
         );
  EDFFX1 \RAM_reg<54><4>  ( .D(n18456), .E(n18349), .CK(clk), .Q(\RAM<54><4> )
         );
  EDFFX1 \RAM_reg<54><3>  ( .D(n18452), .E(n18348), .CK(clk), .Q(\RAM<54><3> )
         );
  EDFFX1 \RAM_reg<54><2>  ( .D(n18448), .E(n18349), .CK(clk), .Q(\RAM<54><2> )
         );
  EDFFX1 \RAM_reg<54><1>  ( .D(n18444), .E(n18348), .CK(clk), .Q(\RAM<54><1> )
         );
  EDFFX1 \RAM_reg<54><0>  ( .D(n18440), .E(n18349), .CK(clk), .Q(\RAM<54><0> )
         );
  EDFFX1 \RAM_reg<46><31>  ( .D(n18564), .E(n18417), .CK(clk), .Q(
        \RAM<46><31> ) );
  EDFFX1 \RAM_reg<46><30>  ( .D(n18560), .E(n18417), .CK(clk), .Q(
        \RAM<46><30> ) );
  EDFFX1 \RAM_reg<46><29>  ( .D(n18556), .E(n18417), .CK(clk), .Q(
        \RAM<46><29> ) );
  EDFFX1 \RAM_reg<46><28>  ( .D(n18552), .E(n18417), .CK(clk), .Q(
        \RAM<46><28> ) );
  EDFFX1 \RAM_reg<46><27>  ( .D(n18548), .E(n18417), .CK(clk), .Q(
        \RAM<46><27> ) );
  EDFFX1 \RAM_reg<46><26>  ( .D(n18544), .E(n18417), .CK(clk), .Q(
        \RAM<46><26> ) );
  EDFFX1 \RAM_reg<46><25>  ( .D(n18540), .E(n18417), .CK(clk), .Q(
        \RAM<46><25> ) );
  EDFFX1 \RAM_reg<46><24>  ( .D(n18536), .E(n18417), .CK(clk), .Q(
        \RAM<46><24> ) );
  EDFFX1 \RAM_reg<46><23>  ( .D(n18532), .E(n18417), .CK(clk), .Q(
        \RAM<46><23> ) );
  EDFFX1 \RAM_reg<46><22>  ( .D(n18528), .E(n18417), .CK(clk), .Q(
        \RAM<46><22> ) );
  EDFFX1 \RAM_reg<46><21>  ( .D(n18524), .E(n18417), .CK(clk), .Q(
        \RAM<46><21> ) );
  EDFFX1 \RAM_reg<46><20>  ( .D(n18520), .E(n18417), .CK(clk), .Q(
        \RAM<46><20> ) );
  EDFFX1 \RAM_reg<46><19>  ( .D(n18516), .E(n18418), .CK(clk), .Q(
        \RAM<46><19> ) );
  EDFFX1 \RAM_reg<46><18>  ( .D(n18512), .E(n18418), .CK(clk), .Q(
        \RAM<46><18> ) );
  EDFFX1 \RAM_reg<46><17>  ( .D(n18508), .E(n18418), .CK(clk), .Q(
        \RAM<46><17> ) );
  EDFFX1 \RAM_reg<46><16>  ( .D(n18504), .E(n18418), .CK(clk), .Q(
        \RAM<46><16> ) );
  EDFFX1 \RAM_reg<46><15>  ( .D(n18500), .E(n18418), .CK(clk), .Q(
        \RAM<46><15> ) );
  EDFFX1 \RAM_reg<46><14>  ( .D(n18496), .E(n18418), .CK(clk), .Q(
        \RAM<46><14> ) );
  EDFFX1 \RAM_reg<46><13>  ( .D(n18492), .E(n18418), .CK(clk), .Q(
        \RAM<46><13> ) );
  EDFFX1 \RAM_reg<46><12>  ( .D(n18488), .E(n18418), .CK(clk), .Q(
        \RAM<46><12> ) );
  EDFFX1 \RAM_reg<46><11>  ( .D(n18484), .E(n18418), .CK(clk), .Q(
        \RAM<46><11> ) );
  EDFFX1 \RAM_reg<46><10>  ( .D(n18480), .E(n18418), .CK(clk), .Q(
        \RAM<46><10> ) );
  EDFFX1 \RAM_reg<46><9>  ( .D(n18476), .E(n18418), .CK(clk), .Q(\RAM<46><9> )
         );
  EDFFX1 \RAM_reg<46><8>  ( .D(n18472), .E(n18418), .CK(clk), .Q(\RAM<46><8> )
         );
  EDFFX1 \RAM_reg<46><7>  ( .D(n18468), .E(n3524), .CK(clk), .Q(\RAM<46><7> )
         );
  EDFFX1 \RAM_reg<46><6>  ( .D(n18464), .E(n3524), .CK(clk), .Q(\RAM<46><6> )
         );
  EDFFX1 \RAM_reg<46><5>  ( .D(n18460), .E(n18417), .CK(clk), .Q(\RAM<46><5> )
         );
  EDFFX1 \RAM_reg<46><4>  ( .D(n18456), .E(n18418), .CK(clk), .Q(\RAM<46><4> )
         );
  EDFFX1 \RAM_reg<46><3>  ( .D(n18452), .E(n18417), .CK(clk), .Q(\RAM<46><3> )
         );
  EDFFX1 \RAM_reg<46><2>  ( .D(n18448), .E(n18418), .CK(clk), .Q(\RAM<46><2> )
         );
  EDFFX1 \RAM_reg<46><1>  ( .D(n18444), .E(n18417), .CK(clk), .Q(\RAM<46><1> )
         );
  EDFFX1 \RAM_reg<46><0>  ( .D(n18440), .E(n18418), .CK(clk), .Q(\RAM<46><0> )
         );
  EDFFX1 \RAM_reg<38><31>  ( .D(n18564), .E(n18411), .CK(clk), .Q(
        \RAM<38><31> ) );
  EDFFX1 \RAM_reg<38><30>  ( .D(n18560), .E(n18411), .CK(clk), .Q(
        \RAM<38><30> ) );
  EDFFX1 \RAM_reg<38><29>  ( .D(n18556), .E(n18411), .CK(clk), .Q(
        \RAM<38><29> ) );
  EDFFX1 \RAM_reg<38><28>  ( .D(n18552), .E(n18411), .CK(clk), .Q(
        \RAM<38><28> ) );
  EDFFX1 \RAM_reg<38><27>  ( .D(n18548), .E(n18411), .CK(clk), .Q(
        \RAM<38><27> ) );
  EDFFX1 \RAM_reg<38><26>  ( .D(n18544), .E(n18411), .CK(clk), .Q(
        \RAM<38><26> ) );
  EDFFX1 \RAM_reg<38><25>  ( .D(n18540), .E(n18411), .CK(clk), .Q(
        \RAM<38><25> ) );
  EDFFX1 \RAM_reg<38><24>  ( .D(n18536), .E(n18411), .CK(clk), .Q(
        \RAM<38><24> ) );
  EDFFX1 \RAM_reg<38><23>  ( .D(n18532), .E(n18411), .CK(clk), .Q(
        \RAM<38><23> ) );
  EDFFX1 \RAM_reg<38><22>  ( .D(n18528), .E(n18411), .CK(clk), .Q(
        \RAM<38><22> ) );
  EDFFX1 \RAM_reg<38><21>  ( .D(n18524), .E(n18411), .CK(clk), .Q(
        \RAM<38><21> ) );
  EDFFX1 \RAM_reg<38><20>  ( .D(n18520), .E(n18411), .CK(clk), .Q(
        \RAM<38><20> ) );
  EDFFX1 \RAM_reg<38><19>  ( .D(n18516), .E(n18412), .CK(clk), .Q(
        \RAM<38><19> ) );
  EDFFX1 \RAM_reg<38><18>  ( .D(n18512), .E(n18412), .CK(clk), .Q(
        \RAM<38><18> ) );
  EDFFX1 \RAM_reg<38><17>  ( .D(n18508), .E(n18412), .CK(clk), .Q(
        \RAM<38><17> ) );
  EDFFX1 \RAM_reg<38><16>  ( .D(n18504), .E(n18412), .CK(clk), .Q(
        \RAM<38><16> ) );
  EDFFX1 \RAM_reg<38><15>  ( .D(n18500), .E(n18412), .CK(clk), .Q(
        \RAM<38><15> ) );
  EDFFX1 \RAM_reg<38><14>  ( .D(n18496), .E(n18412), .CK(clk), .Q(
        \RAM<38><14> ) );
  EDFFX1 \RAM_reg<38><13>  ( .D(n18492), .E(n18412), .CK(clk), .Q(
        \RAM<38><13> ) );
  EDFFX1 \RAM_reg<38><12>  ( .D(n18488), .E(n18412), .CK(clk), .Q(
        \RAM<38><12> ) );
  EDFFX1 \RAM_reg<38><11>  ( .D(n18484), .E(n18412), .CK(clk), .Q(
        \RAM<38><11> ) );
  EDFFX1 \RAM_reg<38><10>  ( .D(n18480), .E(n18412), .CK(clk), .Q(
        \RAM<38><10> ) );
  EDFFX1 \RAM_reg<38><9>  ( .D(n18476), .E(n18412), .CK(clk), .Q(\RAM<38><9> )
         );
  EDFFX1 \RAM_reg<38><8>  ( .D(n18472), .E(n18412), .CK(clk), .Q(\RAM<38><8> )
         );
  EDFFX1 \RAM_reg<38><7>  ( .D(n18468), .E(n3526), .CK(clk), .Q(\RAM<38><7> )
         );
  EDFFX1 \RAM_reg<38><6>  ( .D(n18464), .E(n3526), .CK(clk), .Q(\RAM<38><6> )
         );
  EDFFX1 \RAM_reg<38><5>  ( .D(n18460), .E(n18411), .CK(clk), .Q(\RAM<38><5> )
         );
  EDFFX1 \RAM_reg<38><4>  ( .D(n18456), .E(n18412), .CK(clk), .Q(\RAM<38><4> )
         );
  EDFFX1 \RAM_reg<38><3>  ( .D(n18452), .E(n18411), .CK(clk), .Q(\RAM<38><3> )
         );
  EDFFX1 \RAM_reg<38><2>  ( .D(n18448), .E(n18412), .CK(clk), .Q(\RAM<38><2> )
         );
  EDFFX1 \RAM_reg<38><1>  ( .D(n18444), .E(n18411), .CK(clk), .Q(\RAM<38><1> )
         );
  EDFFX1 \RAM_reg<38><0>  ( .D(n18440), .E(n18412), .CK(clk), .Q(\RAM<38><0> )
         );
  EDFFX1 \RAM_reg<30><31>  ( .D(n18562), .E(n18246), .CK(clk), .Q(
        \RAM<30><31> ) );
  EDFFX1 \RAM_reg<30><30>  ( .D(n18558), .E(n18246), .CK(clk), .Q(
        \RAM<30><30> ) );
  EDFFX1 \RAM_reg<30><29>  ( .D(n18554), .E(n18246), .CK(clk), .Q(
        \RAM<30><29> ) );
  EDFFX1 \RAM_reg<30><28>  ( .D(n18550), .E(n18246), .CK(clk), .Q(
        \RAM<30><28> ) );
  EDFFX1 \RAM_reg<30><27>  ( .D(n18546), .E(n18246), .CK(clk), .Q(
        \RAM<30><27> ) );
  EDFFX1 \RAM_reg<30><26>  ( .D(n18542), .E(n18246), .CK(clk), .Q(
        \RAM<30><26> ) );
  EDFFX1 \RAM_reg<30><25>  ( .D(n18538), .E(n18246), .CK(clk), .Q(
        \RAM<30><25> ) );
  EDFFX1 \RAM_reg<30><24>  ( .D(n18534), .E(n18246), .CK(clk), .Q(
        \RAM<30><24> ) );
  EDFFX1 \RAM_reg<30><23>  ( .D(n18530), .E(n18246), .CK(clk), .Q(
        \RAM<30><23> ) );
  EDFFX1 \RAM_reg<30><22>  ( .D(n18526), .E(n18246), .CK(clk), .Q(
        \RAM<30><22> ) );
  EDFFX1 \RAM_reg<30><21>  ( .D(n18522), .E(n18246), .CK(clk), .Q(
        \RAM<30><21> ) );
  EDFFX1 \RAM_reg<30><20>  ( .D(n18518), .E(n18246), .CK(clk), .Q(
        \RAM<30><20> ) );
  EDFFX1 \RAM_reg<30><19>  ( .D(n18514), .E(n18247), .CK(clk), .Q(
        \RAM<30><19> ) );
  EDFFX1 \RAM_reg<30><18>  ( .D(n18510), .E(n18247), .CK(clk), .Q(
        \RAM<30><18> ) );
  EDFFX1 \RAM_reg<30><17>  ( .D(n18506), .E(n18247), .CK(clk), .Q(
        \RAM<30><17> ) );
  EDFFX1 \RAM_reg<30><16>  ( .D(n18502), .E(n18247), .CK(clk), .Q(
        \RAM<30><16> ) );
  EDFFX1 \RAM_reg<30><15>  ( .D(n18498), .E(n18247), .CK(clk), .Q(
        \RAM<30><15> ) );
  EDFFX1 \RAM_reg<30><14>  ( .D(n18494), .E(n18247), .CK(clk), .Q(
        \RAM<30><14> ) );
  EDFFX1 \RAM_reg<30><13>  ( .D(n18490), .E(n18247), .CK(clk), .Q(
        \RAM<30><13> ) );
  EDFFX1 \RAM_reg<30><12>  ( .D(n18486), .E(n18247), .CK(clk), .Q(
        \RAM<30><12> ) );
  EDFFX1 \RAM_reg<30><11>  ( .D(n18482), .E(n18247), .CK(clk), .Q(
        \RAM<30><11> ) );
  EDFFX1 \RAM_reg<30><10>  ( .D(n18478), .E(n18247), .CK(clk), .Q(
        \RAM<30><10> ) );
  EDFFX1 \RAM_reg<30><9>  ( .D(n18474), .E(n18247), .CK(clk), .Q(\RAM<30><9> )
         );
  EDFFX1 \RAM_reg<30><8>  ( .D(n18470), .E(n18247), .CK(clk), .Q(\RAM<30><8> )
         );
  EDFFX1 \RAM_reg<30><7>  ( .D(n18466), .E(n3576), .CK(clk), .Q(\RAM<30><7> )
         );
  EDFFX1 \RAM_reg<30><6>  ( .D(n18462), .E(n3576), .CK(clk), .Q(\RAM<30><6> )
         );
  EDFFX1 \RAM_reg<30><5>  ( .D(n18458), .E(n18246), .CK(clk), .Q(\RAM<30><5> )
         );
  EDFFX1 \RAM_reg<30><4>  ( .D(n18454), .E(n18247), .CK(clk), .Q(\RAM<30><4> )
         );
  EDFFX1 \RAM_reg<30><3>  ( .D(n18450), .E(n18246), .CK(clk), .Q(\RAM<30><3> )
         );
  EDFFX1 \RAM_reg<30><2>  ( .D(n18446), .E(n18247), .CK(clk), .Q(\RAM<30><2> )
         );
  EDFFX1 \RAM_reg<30><1>  ( .D(n18442), .E(n18246), .CK(clk), .Q(\RAM<30><1> )
         );
  EDFFX1 \RAM_reg<30><0>  ( .D(n18438), .E(n18247), .CK(clk), .Q(\RAM<30><0> )
         );
  EDFFX1 \RAM_reg<22><31>  ( .D(n18564), .E(n18249), .CK(clk), .Q(
        \RAM<22><31> ) );
  EDFFX1 \RAM_reg<22><30>  ( .D(n18560), .E(n18249), .CK(clk), .Q(
        \RAM<22><30> ) );
  EDFFX1 \RAM_reg<22><29>  ( .D(n18556), .E(n18249), .CK(clk), .Q(
        \RAM<22><29> ) );
  EDFFX1 \RAM_reg<22><28>  ( .D(n18552), .E(n18249), .CK(clk), .Q(
        \RAM<22><28> ) );
  EDFFX1 \RAM_reg<22><27>  ( .D(n18548), .E(n18249), .CK(clk), .Q(
        \RAM<22><27> ) );
  EDFFX1 \RAM_reg<22><26>  ( .D(n18544), .E(n18249), .CK(clk), .Q(
        \RAM<22><26> ) );
  EDFFX1 \RAM_reg<22><25>  ( .D(n18540), .E(n18249), .CK(clk), .Q(
        \RAM<22><25> ) );
  EDFFX1 \RAM_reg<22><24>  ( .D(n18536), .E(n18249), .CK(clk), .Q(
        \RAM<22><24> ) );
  EDFFX1 \RAM_reg<22><23>  ( .D(n18532), .E(n18249), .CK(clk), .Q(
        \RAM<22><23> ) );
  EDFFX1 \RAM_reg<22><22>  ( .D(n18528), .E(n18249), .CK(clk), .Q(
        \RAM<22><22> ) );
  EDFFX1 \RAM_reg<22><21>  ( .D(n18524), .E(n18249), .CK(clk), .Q(
        \RAM<22><21> ) );
  EDFFX1 \RAM_reg<22><20>  ( .D(n18520), .E(n18249), .CK(clk), .Q(
        \RAM<22><20> ) );
  EDFFX1 \RAM_reg<22><19>  ( .D(n18516), .E(n18250), .CK(clk), .Q(
        \RAM<22><19> ) );
  EDFFX1 \RAM_reg<22><18>  ( .D(n18512), .E(n18250), .CK(clk), .Q(
        \RAM<22><18> ) );
  EDFFX1 \RAM_reg<22><17>  ( .D(n18508), .E(n18250), .CK(clk), .Q(
        \RAM<22><17> ) );
  EDFFX1 \RAM_reg<22><16>  ( .D(n18504), .E(n18250), .CK(clk), .Q(
        \RAM<22><16> ) );
  EDFFX1 \RAM_reg<22><15>  ( .D(n18500), .E(n18250), .CK(clk), .Q(
        \RAM<22><15> ) );
  EDFFX1 \RAM_reg<22><14>  ( .D(n18496), .E(n18250), .CK(clk), .Q(
        \RAM<22><14> ) );
  EDFFX1 \RAM_reg<22><13>  ( .D(n18492), .E(n18250), .CK(clk), .Q(
        \RAM<22><13> ) );
  EDFFX1 \RAM_reg<22><12>  ( .D(n18488), .E(n18250), .CK(clk), .Q(
        \RAM<22><12> ) );
  EDFFX1 \RAM_reg<22><11>  ( .D(n18484), .E(n18250), .CK(clk), .Q(
        \RAM<22><11> ) );
  EDFFX1 \RAM_reg<22><10>  ( .D(n18480), .E(n18250), .CK(clk), .Q(
        \RAM<22><10> ) );
  EDFFX1 \RAM_reg<22><9>  ( .D(n18476), .E(n18250), .CK(clk), .Q(\RAM<22><9> )
         );
  EDFFX1 \RAM_reg<22><8>  ( .D(n18472), .E(n18250), .CK(clk), .Q(\RAM<22><8> )
         );
  EDFFX1 \RAM_reg<22><7>  ( .D(n18468), .E(n3566), .CK(clk), .Q(\RAM<22><7> )
         );
  EDFFX1 \RAM_reg<22><6>  ( .D(n18464), .E(n3566), .CK(clk), .Q(\RAM<22><6> )
         );
  EDFFX1 \RAM_reg<22><5>  ( .D(n18460), .E(n18249), .CK(clk), .Q(\RAM<22><5> )
         );
  EDFFX1 \RAM_reg<22><4>  ( .D(n18456), .E(n18250), .CK(clk), .Q(\RAM<22><4> )
         );
  EDFFX1 \RAM_reg<22><3>  ( .D(n18452), .E(n18249), .CK(clk), .Q(\RAM<22><3> )
         );
  EDFFX1 \RAM_reg<22><2>  ( .D(n18448), .E(n18250), .CK(clk), .Q(\RAM<22><2> )
         );
  EDFFX1 \RAM_reg<22><1>  ( .D(n18444), .E(n18249), .CK(clk), .Q(\RAM<22><1> )
         );
  EDFFX1 \RAM_reg<22><0>  ( .D(n18440), .E(n18250), .CK(clk), .Q(\RAM<22><0> )
         );
  EDFFX1 \RAM_reg<14><31>  ( .D(n18562), .E(n18252), .CK(clk), .Q(
        \RAM<14><31> ) );
  EDFFX1 \RAM_reg<14><30>  ( .D(n18558), .E(n18252), .CK(clk), .Q(
        \RAM<14><30> ) );
  EDFFX1 \RAM_reg<14><29>  ( .D(n18554), .E(n18252), .CK(clk), .Q(
        \RAM<14><29> ) );
  EDFFX1 \RAM_reg<14><28>  ( .D(n18550), .E(n18252), .CK(clk), .Q(
        \RAM<14><28> ) );
  EDFFX1 \RAM_reg<14><27>  ( .D(n18546), .E(n18252), .CK(clk), .Q(
        \RAM<14><27> ) );
  EDFFX1 \RAM_reg<14><26>  ( .D(n18542), .E(n18252), .CK(clk), .Q(
        \RAM<14><26> ) );
  EDFFX1 \RAM_reg<14><25>  ( .D(n18538), .E(n18252), .CK(clk), .Q(
        \RAM<14><25> ) );
  EDFFX1 \RAM_reg<14><24>  ( .D(n18534), .E(n18252), .CK(clk), .Q(
        \RAM<14><24> ) );
  EDFFX1 \RAM_reg<14><23>  ( .D(n18530), .E(n18252), .CK(clk), .Q(
        \RAM<14><23> ) );
  EDFFX1 \RAM_reg<14><22>  ( .D(n18526), .E(n18252), .CK(clk), .Q(
        \RAM<14><22> ) );
  EDFFX1 \RAM_reg<14><21>  ( .D(n18522), .E(n18252), .CK(clk), .Q(
        \RAM<14><21> ) );
  EDFFX1 \RAM_reg<14><20>  ( .D(n18518), .E(n18252), .CK(clk), .Q(
        \RAM<14><20> ) );
  EDFFX1 \RAM_reg<14><19>  ( .D(n18514), .E(n18253), .CK(clk), .Q(
        \RAM<14><19> ) );
  EDFFX1 \RAM_reg<14><18>  ( .D(n18510), .E(n18253), .CK(clk), .Q(
        \RAM<14><18> ) );
  EDFFX1 \RAM_reg<14><17>  ( .D(n18506), .E(n18253), .CK(clk), .Q(
        \RAM<14><17> ) );
  EDFFX1 \RAM_reg<14><16>  ( .D(n18502), .E(n18253), .CK(clk), .Q(
        \RAM<14><16> ) );
  EDFFX1 \RAM_reg<14><15>  ( .D(n18498), .E(n18253), .CK(clk), .Q(
        \RAM<14><15> ) );
  EDFFX1 \RAM_reg<14><14>  ( .D(n18494), .E(n18253), .CK(clk), .Q(
        \RAM<14><14> ) );
  EDFFX1 \RAM_reg<14><13>  ( .D(n18490), .E(n18253), .CK(clk), .Q(
        \RAM<14><13> ) );
  EDFFX1 \RAM_reg<14><12>  ( .D(n18486), .E(n18253), .CK(clk), .Q(
        \RAM<14><12> ) );
  EDFFX1 \RAM_reg<14><11>  ( .D(n18482), .E(n18253), .CK(clk), .Q(
        \RAM<14><11> ) );
  EDFFX1 \RAM_reg<14><10>  ( .D(n18478), .E(n18253), .CK(clk), .Q(
        \RAM<14><10> ) );
  EDFFX1 \RAM_reg<14><9>  ( .D(n18474), .E(n18253), .CK(clk), .Q(\RAM<14><9> )
         );
  EDFFX1 \RAM_reg<14><8>  ( .D(n18470), .E(n18253), .CK(clk), .Q(\RAM<14><8> )
         );
  EDFFX1 \RAM_reg<14><7>  ( .D(n18466), .E(n3561), .CK(clk), .Q(\RAM<14><7> )
         );
  EDFFX1 \RAM_reg<14><6>  ( .D(n18462), .E(n3561), .CK(clk), .Q(\RAM<14><6> )
         );
  EDFFX1 \RAM_reg<14><5>  ( .D(n18458), .E(n18252), .CK(clk), .Q(\RAM<14><5> )
         );
  EDFFX1 \RAM_reg<14><4>  ( .D(n18454), .E(n18253), .CK(clk), .Q(\RAM<14><4> )
         );
  EDFFX1 \RAM_reg<14><3>  ( .D(n18450), .E(n18252), .CK(clk), .Q(\RAM<14><3> )
         );
  EDFFX1 \RAM_reg<14><2>  ( .D(n18446), .E(n18253), .CK(clk), .Q(\RAM<14><2> )
         );
  EDFFX1 \RAM_reg<14><1>  ( .D(n18442), .E(n18252), .CK(clk), .Q(\RAM<14><1> )
         );
  EDFFX1 \RAM_reg<14><0>  ( .D(n18438), .E(n18253), .CK(clk), .Q(\RAM<14><0> )
         );
  EDFFX1 \RAM_reg<6><31>  ( .D(n18563), .E(n18255), .CK(clk), .Q(\RAM<6><31> )
         );
  EDFFX1 \RAM_reg<6><30>  ( .D(n18559), .E(n18255), .CK(clk), .Q(\RAM<6><30> )
         );
  EDFFX1 \RAM_reg<6><29>  ( .D(n18555), .E(n18255), .CK(clk), .Q(\RAM<6><29> )
         );
  EDFFX1 \RAM_reg<6><28>  ( .D(n18551), .E(n18255), .CK(clk), .Q(\RAM<6><28> )
         );
  EDFFX1 \RAM_reg<6><27>  ( .D(n18547), .E(n18255), .CK(clk), .Q(\RAM<6><27> )
         );
  EDFFX1 \RAM_reg<6><26>  ( .D(n18543), .E(n18255), .CK(clk), .Q(\RAM<6><26> )
         );
  EDFFX1 \RAM_reg<6><25>  ( .D(n18539), .E(n18255), .CK(clk), .Q(\RAM<6><25> )
         );
  EDFFX1 \RAM_reg<6><24>  ( .D(n18535), .E(n18255), .CK(clk), .Q(\RAM<6><24> )
         );
  EDFFX1 \RAM_reg<6><23>  ( .D(n18531), .E(n18255), .CK(clk), .Q(\RAM<6><23> )
         );
  EDFFX1 \RAM_reg<6><22>  ( .D(n18527), .E(n18255), .CK(clk), .Q(\RAM<6><22> )
         );
  EDFFX1 \RAM_reg<6><21>  ( .D(n18523), .E(n18255), .CK(clk), .Q(\RAM<6><21> )
         );
  EDFFX1 \RAM_reg<6><20>  ( .D(n18519), .E(n18255), .CK(clk), .Q(\RAM<6><20> )
         );
  EDFFX1 \RAM_reg<6><19>  ( .D(n18515), .E(n18256), .CK(clk), .Q(\RAM<6><19> )
         );
  EDFFX1 \RAM_reg<6><18>  ( .D(n18511), .E(n18256), .CK(clk), .Q(\RAM<6><18> )
         );
  EDFFX1 \RAM_reg<6><17>  ( .D(n18507), .E(n18256), .CK(clk), .Q(\RAM<6><17> )
         );
  EDFFX1 \RAM_reg<6><16>  ( .D(n18503), .E(n18256), .CK(clk), .Q(\RAM<6><16> )
         );
  EDFFX1 \RAM_reg<6><15>  ( .D(n18499), .E(n18256), .CK(clk), .Q(\RAM<6><15> )
         );
  EDFFX1 \RAM_reg<6><14>  ( .D(n18495), .E(n18256), .CK(clk), .Q(\RAM<6><14> )
         );
  EDFFX1 \RAM_reg<6><13>  ( .D(n18491), .E(n18256), .CK(clk), .Q(\RAM<6><13> )
         );
  EDFFX1 \RAM_reg<6><12>  ( .D(n18487), .E(n18256), .CK(clk), .Q(\RAM<6><12> )
         );
  EDFFX1 \RAM_reg<6><11>  ( .D(n18483), .E(n18256), .CK(clk), .Q(\RAM<6><11> )
         );
  EDFFX1 \RAM_reg<6><10>  ( .D(n18479), .E(n18256), .CK(clk), .Q(\RAM<6><10> )
         );
  EDFFX1 \RAM_reg<6><9>  ( .D(n18475), .E(n18256), .CK(clk), .Q(\RAM<6><9> )
         );
  EDFFX1 \RAM_reg<6><8>  ( .D(n18471), .E(n18256), .CK(clk), .Q(\RAM<6><8> )
         );
  EDFFX1 \RAM_reg<6><7>  ( .D(n18467), .E(n3560), .CK(clk), .Q(\RAM<6><7> ) );
  EDFFX1 \RAM_reg<6><6>  ( .D(n18463), .E(n3560), .CK(clk), .Q(\RAM<6><6> ) );
  EDFFX1 \RAM_reg<6><5>  ( .D(n18459), .E(n18255), .CK(clk), .Q(\RAM<6><5> )
         );
  EDFFX1 \RAM_reg<6><4>  ( .D(n18455), .E(n18256), .CK(clk), .Q(\RAM<6><4> )
         );
  EDFFX1 \RAM_reg<6><3>  ( .D(n18451), .E(n18255), .CK(clk), .Q(\RAM<6><3> )
         );
  EDFFX1 \RAM_reg<6><2>  ( .D(n18447), .E(n18256), .CK(clk), .Q(\RAM<6><2> )
         );
  EDFFX1 \RAM_reg<6><1>  ( .D(n18443), .E(n18255), .CK(clk), .Q(\RAM<6><1> )
         );
  EDFFX1 \RAM_reg<6><0>  ( .D(n18439), .E(n18256), .CK(clk), .Q(\RAM<6><0> )
         );
  EDFFX1 \RAM_reg<61><31>  ( .D(n18562), .E(n18363), .CK(clk), .Q(
        \RAM<61><31> ) );
  EDFFX1 \RAM_reg<61><30>  ( .D(n18558), .E(n18363), .CK(clk), .Q(
        \RAM<61><30> ) );
  EDFFX1 \RAM_reg<61><29>  ( .D(n18554), .E(n18363), .CK(clk), .Q(
        \RAM<61><29> ) );
  EDFFX1 \RAM_reg<61><28>  ( .D(n18550), .E(n18363), .CK(clk), .Q(
        \RAM<61><28> ) );
  EDFFX1 \RAM_reg<61><27>  ( .D(n18546), .E(n18363), .CK(clk), .Q(
        \RAM<61><27> ) );
  EDFFX1 \RAM_reg<61><26>  ( .D(n18542), .E(n18363), .CK(clk), .Q(
        \RAM<61><26> ) );
  EDFFX1 \RAM_reg<61><25>  ( .D(n18538), .E(n18363), .CK(clk), .Q(
        \RAM<61><25> ) );
  EDFFX1 \RAM_reg<61><24>  ( .D(n18534), .E(n18363), .CK(clk), .Q(
        \RAM<61><24> ) );
  EDFFX1 \RAM_reg<61><23>  ( .D(n18530), .E(n18363), .CK(clk), .Q(
        \RAM<61><23> ) );
  EDFFX1 \RAM_reg<61><22>  ( .D(n18526), .E(n18363), .CK(clk), .Q(
        \RAM<61><22> ) );
  EDFFX1 \RAM_reg<61><21>  ( .D(n18522), .E(n18363), .CK(clk), .Q(
        \RAM<61><21> ) );
  EDFFX1 \RAM_reg<61><20>  ( .D(n18518), .E(n18363), .CK(clk), .Q(
        \RAM<61><20> ) );
  EDFFX1 \RAM_reg<61><19>  ( .D(n18514), .E(n18364), .CK(clk), .Q(
        \RAM<61><19> ) );
  EDFFX1 \RAM_reg<61><18>  ( .D(n18510), .E(n18364), .CK(clk), .Q(
        \RAM<61><18> ) );
  EDFFX1 \RAM_reg<61><17>  ( .D(n18506), .E(n18364), .CK(clk), .Q(
        \RAM<61><17> ) );
  EDFFX1 \RAM_reg<61><16>  ( .D(n18502), .E(n18364), .CK(clk), .Q(
        \RAM<61><16> ) );
  EDFFX1 \RAM_reg<61><15>  ( .D(n18498), .E(n18364), .CK(clk), .Q(
        \RAM<61><15> ) );
  EDFFX1 \RAM_reg<61><14>  ( .D(n18494), .E(n18364), .CK(clk), .Q(
        \RAM<61><14> ) );
  EDFFX1 \RAM_reg<61><13>  ( .D(n18490), .E(n18364), .CK(clk), .Q(
        \RAM<61><13> ) );
  EDFFX1 \RAM_reg<61><12>  ( .D(n18486), .E(n18364), .CK(clk), .Q(
        \RAM<61><12> ) );
  EDFFX1 \RAM_reg<61><11>  ( .D(n18482), .E(n18364), .CK(clk), .Q(
        \RAM<61><11> ) );
  EDFFX1 \RAM_reg<61><10>  ( .D(n18478), .E(n18364), .CK(clk), .Q(
        \RAM<61><10> ) );
  EDFFX1 \RAM_reg<61><9>  ( .D(n18474), .E(n18364), .CK(clk), .Q(\RAM<61><9> )
         );
  EDFFX1 \RAM_reg<61><8>  ( .D(n18470), .E(n18364), .CK(clk), .Q(\RAM<61><8> )
         );
  EDFFX1 \RAM_reg<61><7>  ( .D(n18466), .E(n3543), .CK(clk), .Q(\RAM<61><7> )
         );
  EDFFX1 \RAM_reg<61><6>  ( .D(n18462), .E(n3543), .CK(clk), .Q(\RAM<61><6> )
         );
  EDFFX1 \RAM_reg<61><5>  ( .D(n18458), .E(n18363), .CK(clk), .Q(\RAM<61><5> )
         );
  EDFFX1 \RAM_reg<61><4>  ( .D(n18454), .E(n18364), .CK(clk), .Q(\RAM<61><4> )
         );
  EDFFX1 \RAM_reg<61><3>  ( .D(n18450), .E(n18363), .CK(clk), .Q(\RAM<61><3> )
         );
  EDFFX1 \RAM_reg<61><2>  ( .D(n18446), .E(n18364), .CK(clk), .Q(\RAM<61><2> )
         );
  EDFFX1 \RAM_reg<61><1>  ( .D(n18442), .E(n18363), .CK(clk), .Q(\RAM<61><1> )
         );
  EDFFX1 \RAM_reg<61><0>  ( .D(n18438), .E(n18364), .CK(clk), .Q(\RAM<61><0> )
         );
  EDFFX1 \RAM_reg<53><31>  ( .D(n18562), .E(n18345), .CK(clk), .Q(
        \RAM<53><31> ) );
  EDFFX1 \RAM_reg<53><30>  ( .D(n18558), .E(n18345), .CK(clk), .Q(
        \RAM<53><30> ) );
  EDFFX1 \RAM_reg<53><29>  ( .D(n18554), .E(n18345), .CK(clk), .Q(
        \RAM<53><29> ) );
  EDFFX1 \RAM_reg<53><28>  ( .D(n18550), .E(n18345), .CK(clk), .Q(
        \RAM<53><28> ) );
  EDFFX1 \RAM_reg<53><27>  ( .D(n18546), .E(n18345), .CK(clk), .Q(
        \RAM<53><27> ) );
  EDFFX1 \RAM_reg<53><26>  ( .D(n18542), .E(n18345), .CK(clk), .Q(
        \RAM<53><26> ) );
  EDFFX1 \RAM_reg<53><25>  ( .D(n18538), .E(n18345), .CK(clk), .Q(
        \RAM<53><25> ) );
  EDFFX1 \RAM_reg<53><24>  ( .D(n18534), .E(n18345), .CK(clk), .Q(
        \RAM<53><24> ) );
  EDFFX1 \RAM_reg<53><23>  ( .D(n18530), .E(n18345), .CK(clk), .Q(
        \RAM<53><23> ) );
  EDFFX1 \RAM_reg<53><22>  ( .D(n18526), .E(n18345), .CK(clk), .Q(
        \RAM<53><22> ) );
  EDFFX1 \RAM_reg<53><21>  ( .D(n18522), .E(n18345), .CK(clk), .Q(
        \RAM<53><21> ) );
  EDFFX1 \RAM_reg<53><20>  ( .D(n18518), .E(n18345), .CK(clk), .Q(
        \RAM<53><20> ) );
  EDFFX1 \RAM_reg<53><19>  ( .D(n18514), .E(n18346), .CK(clk), .Q(
        \RAM<53><19> ) );
  EDFFX1 \RAM_reg<53><18>  ( .D(n18510), .E(n18346), .CK(clk), .Q(
        \RAM<53><18> ) );
  EDFFX1 \RAM_reg<53><17>  ( .D(n18506), .E(n18346), .CK(clk), .Q(
        \RAM<53><17> ) );
  EDFFX1 \RAM_reg<53><16>  ( .D(n18502), .E(n18346), .CK(clk), .Q(
        \RAM<53><16> ) );
  EDFFX1 \RAM_reg<53><15>  ( .D(n18498), .E(n18346), .CK(clk), .Q(
        \RAM<53><15> ) );
  EDFFX1 \RAM_reg<53><14>  ( .D(n18494), .E(n18346), .CK(clk), .Q(
        \RAM<53><14> ) );
  EDFFX1 \RAM_reg<53><13>  ( .D(n18490), .E(n18346), .CK(clk), .Q(
        \RAM<53><13> ) );
  EDFFX1 \RAM_reg<53><12>  ( .D(n18486), .E(n18346), .CK(clk), .Q(
        \RAM<53><12> ) );
  EDFFX1 \RAM_reg<53><11>  ( .D(n18482), .E(n18346), .CK(clk), .Q(
        \RAM<53><11> ) );
  EDFFX1 \RAM_reg<53><10>  ( .D(n18478), .E(n18346), .CK(clk), .Q(
        \RAM<53><10> ) );
  EDFFX1 \RAM_reg<53><9>  ( .D(n18474), .E(n18346), .CK(clk), .Q(\RAM<53><9> )
         );
  EDFFX1 \RAM_reg<53><8>  ( .D(n18470), .E(n18346), .CK(clk), .Q(\RAM<53><8> )
         );
  EDFFX1 \RAM_reg<53><7>  ( .D(n18466), .E(n3550), .CK(clk), .Q(\RAM<53><7> )
         );
  EDFFX1 \RAM_reg<53><6>  ( .D(n18462), .E(n3550), .CK(clk), .Q(\RAM<53><6> )
         );
  EDFFX1 \RAM_reg<53><5>  ( .D(n18458), .E(n18345), .CK(clk), .Q(\RAM<53><5> )
         );
  EDFFX1 \RAM_reg<53><4>  ( .D(n18454), .E(n18346), .CK(clk), .Q(\RAM<53><4> )
         );
  EDFFX1 \RAM_reg<53><3>  ( .D(n18450), .E(n18345), .CK(clk), .Q(\RAM<53><3> )
         );
  EDFFX1 \RAM_reg<53><2>  ( .D(n18446), .E(n18346), .CK(clk), .Q(\RAM<53><2> )
         );
  EDFFX1 \RAM_reg<53><1>  ( .D(n18442), .E(n18345), .CK(clk), .Q(\RAM<53><1> )
         );
  EDFFX1 \RAM_reg<53><0>  ( .D(n18438), .E(n18346), .CK(clk), .Q(\RAM<53><0> )
         );
  EDFFX1 \RAM_reg<45><31>  ( .D(n18562), .E(n18375), .CK(clk), .Q(
        \RAM<45><31> ) );
  EDFFX1 \RAM_reg<45><30>  ( .D(n18558), .E(n18375), .CK(clk), .Q(
        \RAM<45><30> ) );
  EDFFX1 \RAM_reg<45><29>  ( .D(n18554), .E(n18375), .CK(clk), .Q(
        \RAM<45><29> ) );
  EDFFX1 \RAM_reg<45><28>  ( .D(n18550), .E(n18375), .CK(clk), .Q(
        \RAM<45><28> ) );
  EDFFX1 \RAM_reg<45><27>  ( .D(n18546), .E(n18375), .CK(clk), .Q(
        \RAM<45><27> ) );
  EDFFX1 \RAM_reg<45><26>  ( .D(n18542), .E(n18375), .CK(clk), .Q(
        \RAM<45><26> ) );
  EDFFX1 \RAM_reg<45><25>  ( .D(n18538), .E(n18375), .CK(clk), .Q(
        \RAM<45><25> ) );
  EDFFX1 \RAM_reg<45><24>  ( .D(n18534), .E(n18375), .CK(clk), .Q(
        \RAM<45><24> ) );
  EDFFX1 \RAM_reg<45><23>  ( .D(n18530), .E(n18375), .CK(clk), .Q(
        \RAM<45><23> ) );
  EDFFX1 \RAM_reg<45><22>  ( .D(n18526), .E(n18375), .CK(clk), .Q(
        \RAM<45><22> ) );
  EDFFX1 \RAM_reg<45><21>  ( .D(n18522), .E(n18375), .CK(clk), .Q(
        \RAM<45><21> ) );
  EDFFX1 \RAM_reg<45><20>  ( .D(n18518), .E(n18375), .CK(clk), .Q(
        \RAM<45><20> ) );
  EDFFX1 \RAM_reg<45><19>  ( .D(n18514), .E(n18376), .CK(clk), .Q(
        \RAM<45><19> ) );
  EDFFX1 \RAM_reg<45><18>  ( .D(n18510), .E(n18376), .CK(clk), .Q(
        \RAM<45><18> ) );
  EDFFX1 \RAM_reg<45><17>  ( .D(n18506), .E(n18376), .CK(clk), .Q(
        \RAM<45><17> ) );
  EDFFX1 \RAM_reg<45><16>  ( .D(n18502), .E(n18376), .CK(clk), .Q(
        \RAM<45><16> ) );
  EDFFX1 \RAM_reg<45><15>  ( .D(n18498), .E(n18376), .CK(clk), .Q(
        \RAM<45><15> ) );
  EDFFX1 \RAM_reg<45><14>  ( .D(n18494), .E(n18376), .CK(clk), .Q(
        \RAM<45><14> ) );
  EDFFX1 \RAM_reg<45><13>  ( .D(n18490), .E(n18376), .CK(clk), .Q(
        \RAM<45><13> ) );
  EDFFX1 \RAM_reg<45><12>  ( .D(n18486), .E(n18376), .CK(clk), .Q(
        \RAM<45><12> ) );
  EDFFX1 \RAM_reg<45><11>  ( .D(n18482), .E(n18376), .CK(clk), .Q(
        \RAM<45><11> ) );
  EDFFX1 \RAM_reg<45><10>  ( .D(n18478), .E(n18376), .CK(clk), .Q(
        \RAM<45><10> ) );
  EDFFX1 \RAM_reg<45><9>  ( .D(n18474), .E(n18376), .CK(clk), .Q(\RAM<45><9> )
         );
  EDFFX1 \RAM_reg<45><8>  ( .D(n18470), .E(n18376), .CK(clk), .Q(\RAM<45><8> )
         );
  EDFFX1 \RAM_reg<45><7>  ( .D(n18466), .E(n3539), .CK(clk), .Q(\RAM<45><7> )
         );
  EDFFX1 \RAM_reg<45><6>  ( .D(n18462), .E(n3539), .CK(clk), .Q(\RAM<45><6> )
         );
  EDFFX1 \RAM_reg<45><5>  ( .D(n18458), .E(n18375), .CK(clk), .Q(\RAM<45><5> )
         );
  EDFFX1 \RAM_reg<45><4>  ( .D(n18454), .E(n18376), .CK(clk), .Q(\RAM<45><4> )
         );
  EDFFX1 \RAM_reg<45><3>  ( .D(n18450), .E(n18375), .CK(clk), .Q(\RAM<45><3> )
         );
  EDFFX1 \RAM_reg<45><2>  ( .D(n18446), .E(n18376), .CK(clk), .Q(\RAM<45><2> )
         );
  EDFFX1 \RAM_reg<45><1>  ( .D(n18442), .E(n18375), .CK(clk), .Q(\RAM<45><1> )
         );
  EDFFX1 \RAM_reg<45><0>  ( .D(n18438), .E(n18376), .CK(clk), .Q(\RAM<45><0> )
         );
  EDFFX1 \RAM_reg<37><31>  ( .D(n18562), .E(n18414), .CK(clk), .Q(
        \RAM<37><31> ) );
  EDFFX1 \RAM_reg<37><30>  ( .D(n18558), .E(n18414), .CK(clk), .Q(
        \RAM<37><30> ) );
  EDFFX1 \RAM_reg<37><29>  ( .D(n18554), .E(n18414), .CK(clk), .Q(
        \RAM<37><29> ) );
  EDFFX1 \RAM_reg<37><28>  ( .D(n18550), .E(n18414), .CK(clk), .Q(
        \RAM<37><28> ) );
  EDFFX1 \RAM_reg<37><27>  ( .D(n18546), .E(n18414), .CK(clk), .Q(
        \RAM<37><27> ) );
  EDFFX1 \RAM_reg<37><26>  ( .D(n18542), .E(n18414), .CK(clk), .Q(
        \RAM<37><26> ) );
  EDFFX1 \RAM_reg<37><25>  ( .D(n18538), .E(n18414), .CK(clk), .Q(
        \RAM<37><25> ) );
  EDFFX1 \RAM_reg<37><24>  ( .D(n18534), .E(n18414), .CK(clk), .Q(
        \RAM<37><24> ) );
  EDFFX1 \RAM_reg<37><23>  ( .D(n18530), .E(n18414), .CK(clk), .Q(
        \RAM<37><23> ) );
  EDFFX1 \RAM_reg<37><22>  ( .D(n18526), .E(n18414), .CK(clk), .Q(
        \RAM<37><22> ) );
  EDFFX1 \RAM_reg<37><21>  ( .D(n18522), .E(n18414), .CK(clk), .Q(
        \RAM<37><21> ) );
  EDFFX1 \RAM_reg<37><20>  ( .D(n18518), .E(n18414), .CK(clk), .Q(
        \RAM<37><20> ) );
  EDFFX1 \RAM_reg<37><19>  ( .D(n18514), .E(n18415), .CK(clk), .Q(
        \RAM<37><19> ) );
  EDFFX1 \RAM_reg<37><18>  ( .D(n18510), .E(n18415), .CK(clk), .Q(
        \RAM<37><18> ) );
  EDFFX1 \RAM_reg<37><17>  ( .D(n18506), .E(n18415), .CK(clk), .Q(
        \RAM<37><17> ) );
  EDFFX1 \RAM_reg<37><16>  ( .D(n18502), .E(n18415), .CK(clk), .Q(
        \RAM<37><16> ) );
  EDFFX1 \RAM_reg<37><15>  ( .D(n18498), .E(n18415), .CK(clk), .Q(
        \RAM<37><15> ) );
  EDFFX1 \RAM_reg<37><14>  ( .D(n18494), .E(n18415), .CK(clk), .Q(
        \RAM<37><14> ) );
  EDFFX1 \RAM_reg<37><13>  ( .D(n18490), .E(n18415), .CK(clk), .Q(
        \RAM<37><13> ) );
  EDFFX1 \RAM_reg<37><12>  ( .D(n18486), .E(n18415), .CK(clk), .Q(
        \RAM<37><12> ) );
  EDFFX1 \RAM_reg<37><11>  ( .D(n18482), .E(n18415), .CK(clk), .Q(
        \RAM<37><11> ) );
  EDFFX1 \RAM_reg<37><10>  ( .D(n18478), .E(n18415), .CK(clk), .Q(
        \RAM<37><10> ) );
  EDFFX1 \RAM_reg<37><9>  ( .D(n18474), .E(n18415), .CK(clk), .Q(\RAM<37><9> )
         );
  EDFFX1 \RAM_reg<37><8>  ( .D(n18470), .E(n18415), .CK(clk), .Q(\RAM<37><8> )
         );
  EDFFX1 \RAM_reg<37><7>  ( .D(n18466), .E(n3525), .CK(clk), .Q(\RAM<37><7> )
         );
  EDFFX1 \RAM_reg<37><6>  ( .D(n18462), .E(n3525), .CK(clk), .Q(\RAM<37><6> )
         );
  EDFFX1 \RAM_reg<37><5>  ( .D(n18458), .E(n18414), .CK(clk), .Q(\RAM<37><5> )
         );
  EDFFX1 \RAM_reg<37><4>  ( .D(n18454), .E(n18415), .CK(clk), .Q(\RAM<37><4> )
         );
  EDFFX1 \RAM_reg<37><3>  ( .D(n18450), .E(n18414), .CK(clk), .Q(\RAM<37><3> )
         );
  EDFFX1 \RAM_reg<37><2>  ( .D(n18446), .E(n18415), .CK(clk), .Q(\RAM<37><2> )
         );
  EDFFX1 \RAM_reg<37><1>  ( .D(n18442), .E(n18414), .CK(clk), .Q(\RAM<37><1> )
         );
  EDFFX1 \RAM_reg<37><0>  ( .D(n18438), .E(n18415), .CK(clk), .Q(\RAM<37><0> )
         );
  EDFFX1 \RAM_reg<29><31>  ( .D(n18562), .E(n18294), .CK(clk), .Q(
        \RAM<29><31> ) );
  EDFFX1 \RAM_reg<29><30>  ( .D(n18558), .E(n18294), .CK(clk), .Q(
        \RAM<29><30> ) );
  EDFFX1 \RAM_reg<29><29>  ( .D(n18554), .E(n18294), .CK(clk), .Q(
        \RAM<29><29> ) );
  EDFFX1 \RAM_reg<29><28>  ( .D(n18550), .E(n18294), .CK(clk), .Q(
        \RAM<29><28> ) );
  EDFFX1 \RAM_reg<29><27>  ( .D(n18546), .E(n18294), .CK(clk), .Q(
        \RAM<29><27> ) );
  EDFFX1 \RAM_reg<29><26>  ( .D(n18542), .E(n18294), .CK(clk), .Q(
        \RAM<29><26> ) );
  EDFFX1 \RAM_reg<29><25>  ( .D(n18538), .E(n18294), .CK(clk), .Q(
        \RAM<29><25> ) );
  EDFFX1 \RAM_reg<29><24>  ( .D(n18534), .E(n18294), .CK(clk), .Q(
        \RAM<29><24> ) );
  EDFFX1 \RAM_reg<29><23>  ( .D(n18530), .E(n18294), .CK(clk), .Q(
        \RAM<29><23> ) );
  EDFFX1 \RAM_reg<29><22>  ( .D(n18526), .E(n18294), .CK(clk), .Q(
        \RAM<29><22> ) );
  EDFFX1 \RAM_reg<29><21>  ( .D(n18522), .E(n18294), .CK(clk), .Q(
        \RAM<29><21> ) );
  EDFFX1 \RAM_reg<29><20>  ( .D(n18518), .E(n18294), .CK(clk), .Q(
        \RAM<29><20> ) );
  EDFFX1 \RAM_reg<29><19>  ( .D(n18514), .E(n18295), .CK(clk), .Q(
        \RAM<29><19> ) );
  EDFFX1 \RAM_reg<29><18>  ( .D(n18510), .E(n18295), .CK(clk), .Q(
        \RAM<29><18> ) );
  EDFFX1 \RAM_reg<29><17>  ( .D(n18506), .E(n18295), .CK(clk), .Q(
        \RAM<29><17> ) );
  EDFFX1 \RAM_reg<29><16>  ( .D(n18502), .E(n18295), .CK(clk), .Q(
        \RAM<29><16> ) );
  EDFFX1 \RAM_reg<29><15>  ( .D(n18498), .E(n18295), .CK(clk), .Q(
        \RAM<29><15> ) );
  EDFFX1 \RAM_reg<29><14>  ( .D(n18494), .E(n18295), .CK(clk), .Q(
        \RAM<29><14> ) );
  EDFFX1 \RAM_reg<29><13>  ( .D(n18490), .E(n18295), .CK(clk), .Q(
        \RAM<29><13> ) );
  EDFFX1 \RAM_reg<29><12>  ( .D(n18486), .E(n18295), .CK(clk), .Q(
        \RAM<29><12> ) );
  EDFFX1 \RAM_reg<29><11>  ( .D(n18482), .E(n18295), .CK(clk), .Q(
        \RAM<29><11> ) );
  EDFFX1 \RAM_reg<29><10>  ( .D(n18478), .E(n18295), .CK(clk), .Q(
        \RAM<29><10> ) );
  EDFFX1 \RAM_reg<29><9>  ( .D(n18474), .E(n18295), .CK(clk), .Q(\RAM<29><9> )
         );
  EDFFX1 \RAM_reg<29><8>  ( .D(n18470), .E(n18295), .CK(clk), .Q(\RAM<29><8> )
         );
  EDFFX1 \RAM_reg<29><7>  ( .D(n18466), .E(n3572), .CK(clk), .Q(\RAM<29><7> )
         );
  EDFFX1 \RAM_reg<29><6>  ( .D(n18462), .E(n3572), .CK(clk), .Q(\RAM<29><6> )
         );
  EDFFX1 \RAM_reg<29><5>  ( .D(n18458), .E(n18294), .CK(clk), .Q(\RAM<29><5> )
         );
  EDFFX1 \RAM_reg<29><4>  ( .D(n18454), .E(n18295), .CK(clk), .Q(\RAM<29><4> )
         );
  EDFFX1 \RAM_reg<29><3>  ( .D(n18450), .E(n18294), .CK(clk), .Q(\RAM<29><3> )
         );
  EDFFX1 \RAM_reg<29><2>  ( .D(n18446), .E(n18295), .CK(clk), .Q(\RAM<29><2> )
         );
  EDFFX1 \RAM_reg<29><1>  ( .D(n18442), .E(n18294), .CK(clk), .Q(\RAM<29><1> )
         );
  EDFFX1 \RAM_reg<29><0>  ( .D(n18438), .E(n18295), .CK(clk), .Q(\RAM<29><0> )
         );
  EDFFX1 \RAM_reg<21><31>  ( .D(n18562), .E(n18369), .CK(clk), .Q(
        \RAM<21><31> ) );
  EDFFX1 \RAM_reg<21><30>  ( .D(n18558), .E(n18369), .CK(clk), .Q(
        \RAM<21><30> ) );
  EDFFX1 \RAM_reg<21><29>  ( .D(n18554), .E(n18369), .CK(clk), .Q(
        \RAM<21><29> ) );
  EDFFX1 \RAM_reg<21><28>  ( .D(n18550), .E(n18369), .CK(clk), .Q(
        \RAM<21><28> ) );
  EDFFX1 \RAM_reg<21><27>  ( .D(n18546), .E(n18369), .CK(clk), .Q(
        \RAM<21><27> ) );
  EDFFX1 \RAM_reg<21><26>  ( .D(n18542), .E(n18369), .CK(clk), .Q(
        \RAM<21><26> ) );
  EDFFX1 \RAM_reg<21><25>  ( .D(n18538), .E(n18369), .CK(clk), .Q(
        \RAM<21><25> ) );
  EDFFX1 \RAM_reg<21><24>  ( .D(n18534), .E(n18369), .CK(clk), .Q(
        \RAM<21><24> ) );
  EDFFX1 \RAM_reg<21><23>  ( .D(n18530), .E(n18369), .CK(clk), .Q(
        \RAM<21><23> ) );
  EDFFX1 \RAM_reg<21><22>  ( .D(n18526), .E(n18369), .CK(clk), .Q(
        \RAM<21><22> ) );
  EDFFX1 \RAM_reg<21><21>  ( .D(n18522), .E(n18369), .CK(clk), .Q(
        \RAM<21><21> ) );
  EDFFX1 \RAM_reg<21><20>  ( .D(n18518), .E(n18369), .CK(clk), .Q(
        \RAM<21><20> ) );
  EDFFX1 \RAM_reg<21><19>  ( .D(n18514), .E(n18370), .CK(clk), .Q(
        \RAM<21><19> ) );
  EDFFX1 \RAM_reg<21><18>  ( .D(n18510), .E(n18370), .CK(clk), .Q(
        \RAM<21><18> ) );
  EDFFX1 \RAM_reg<21><17>  ( .D(n18506), .E(n18370), .CK(clk), .Q(
        \RAM<21><17> ) );
  EDFFX1 \RAM_reg<21><16>  ( .D(n18502), .E(n18370), .CK(clk), .Q(
        \RAM<21><16> ) );
  EDFFX1 \RAM_reg<21><15>  ( .D(n18498), .E(n18370), .CK(clk), .Q(
        \RAM<21><15> ) );
  EDFFX1 \RAM_reg<21><14>  ( .D(n18494), .E(n18370), .CK(clk), .Q(
        \RAM<21><14> ) );
  EDFFX1 \RAM_reg<21><13>  ( .D(n18490), .E(n18370), .CK(clk), .Q(
        \RAM<21><13> ) );
  EDFFX1 \RAM_reg<21><12>  ( .D(n18486), .E(n18370), .CK(clk), .Q(
        \RAM<21><12> ) );
  EDFFX1 \RAM_reg<21><11>  ( .D(n18482), .E(n18370), .CK(clk), .Q(
        \RAM<21><11> ) );
  EDFFX1 \RAM_reg<21><10>  ( .D(n18478), .E(n18370), .CK(clk), .Q(
        \RAM<21><10> ) );
  EDFFX1 \RAM_reg<21><9>  ( .D(n18474), .E(n18370), .CK(clk), .Q(\RAM<21><9> )
         );
  EDFFX1 \RAM_reg<21><8>  ( .D(n18470), .E(n18370), .CK(clk), .Q(\RAM<21><8> )
         );
  EDFFX1 \RAM_reg<21><7>  ( .D(n18466), .E(n3541), .CK(clk), .Q(\RAM<21><7> )
         );
  EDFFX1 \RAM_reg<21><6>  ( .D(n18462), .E(n3541), .CK(clk), .Q(\RAM<21><6> )
         );
  EDFFX1 \RAM_reg<21><5>  ( .D(n18458), .E(n18369), .CK(clk), .Q(\RAM<21><5> )
         );
  EDFFX1 \RAM_reg<21><4>  ( .D(n18454), .E(n18370), .CK(clk), .Q(\RAM<21><4> )
         );
  EDFFX1 \RAM_reg<21><3>  ( .D(n18450), .E(n18369), .CK(clk), .Q(\RAM<21><3> )
         );
  EDFFX1 \RAM_reg<21><2>  ( .D(n18446), .E(n18370), .CK(clk), .Q(\RAM<21><2> )
         );
  EDFFX1 \RAM_reg<21><1>  ( .D(n18442), .E(n18369), .CK(clk), .Q(\RAM<21><1> )
         );
  EDFFX1 \RAM_reg<21><0>  ( .D(n18438), .E(n18370), .CK(clk), .Q(\RAM<21><0> )
         );
  EDFFX1 \RAM_reg<13><31>  ( .D(n18562), .E(n18285), .CK(clk), .Q(
        \RAM<13><31> ) );
  EDFFX1 \RAM_reg<13><30>  ( .D(n18558), .E(n18285), .CK(clk), .Q(
        \RAM<13><30> ) );
  EDFFX1 \RAM_reg<13><29>  ( .D(n18554), .E(n18285), .CK(clk), .Q(
        \RAM<13><29> ) );
  EDFFX1 \RAM_reg<13><28>  ( .D(n18550), .E(n18285), .CK(clk), .Q(
        \RAM<13><28> ) );
  EDFFX1 \RAM_reg<13><27>  ( .D(n18546), .E(n18285), .CK(clk), .Q(
        \RAM<13><27> ) );
  EDFFX1 \RAM_reg<13><26>  ( .D(n18542), .E(n18285), .CK(clk), .Q(
        \RAM<13><26> ) );
  EDFFX1 \RAM_reg<13><25>  ( .D(n18538), .E(n18285), .CK(clk), .Q(
        \RAM<13><25> ) );
  EDFFX1 \RAM_reg<13><24>  ( .D(n18534), .E(n18285), .CK(clk), .Q(
        \RAM<13><24> ) );
  EDFFX1 \RAM_reg<13><23>  ( .D(n18530), .E(n18285), .CK(clk), .Q(
        \RAM<13><23> ) );
  EDFFX1 \RAM_reg<13><22>  ( .D(n18526), .E(n18285), .CK(clk), .Q(
        \RAM<13><22> ) );
  EDFFX1 \RAM_reg<13><21>  ( .D(n18522), .E(n18285), .CK(clk), .Q(
        \RAM<13><21> ) );
  EDFFX1 \RAM_reg<13><20>  ( .D(n18518), .E(n18285), .CK(clk), .Q(
        \RAM<13><20> ) );
  EDFFX1 \RAM_reg<13><19>  ( .D(n18514), .E(n18286), .CK(clk), .Q(
        \RAM<13><19> ) );
  EDFFX1 \RAM_reg<13><18>  ( .D(n18510), .E(n18286), .CK(clk), .Q(
        \RAM<13><18> ) );
  EDFFX1 \RAM_reg<13><17>  ( .D(n18506), .E(n18286), .CK(clk), .Q(
        \RAM<13><17> ) );
  EDFFX1 \RAM_reg<13><16>  ( .D(n18502), .E(n18286), .CK(clk), .Q(
        \RAM<13><16> ) );
  EDFFX1 \RAM_reg<13><15>  ( .D(n18498), .E(n18286), .CK(clk), .Q(
        \RAM<13><15> ) );
  EDFFX1 \RAM_reg<13><14>  ( .D(n18494), .E(n18286), .CK(clk), .Q(
        \RAM<13><14> ) );
  EDFFX1 \RAM_reg<13><13>  ( .D(n18490), .E(n18286), .CK(clk), .Q(
        \RAM<13><13> ) );
  EDFFX1 \RAM_reg<13><12>  ( .D(n18486), .E(n18286), .CK(clk), .Q(
        \RAM<13><12> ) );
  EDFFX1 \RAM_reg<13><11>  ( .D(n18482), .E(n18286), .CK(clk), .Q(
        \RAM<13><11> ) );
  EDFFX1 \RAM_reg<13><10>  ( .D(n18478), .E(n18286), .CK(clk), .Q(
        \RAM<13><10> ) );
  EDFFX1 \RAM_reg<13><9>  ( .D(n18474), .E(n18286), .CK(clk), .Q(\RAM<13><9> )
         );
  EDFFX1 \RAM_reg<13><8>  ( .D(n18470), .E(n18286), .CK(clk), .Q(\RAM<13><8> )
         );
  EDFFX1 \RAM_reg<13><7>  ( .D(n18466), .E(n3575), .CK(clk), .Q(\RAM<13><7> )
         );
  EDFFX1 \RAM_reg<13><6>  ( .D(n18462), .E(n3575), .CK(clk), .Q(\RAM<13><6> )
         );
  EDFFX1 \RAM_reg<13><5>  ( .D(n18458), .E(n18285), .CK(clk), .Q(\RAM<13><5> )
         );
  EDFFX1 \RAM_reg<13><4>  ( .D(n18454), .E(n18286), .CK(clk), .Q(\RAM<13><4> )
         );
  EDFFX1 \RAM_reg<13><3>  ( .D(n18450), .E(n18285), .CK(clk), .Q(\RAM<13><3> )
         );
  EDFFX1 \RAM_reg<13><2>  ( .D(n18446), .E(n18286), .CK(clk), .Q(\RAM<13><2> )
         );
  EDFFX1 \RAM_reg<13><1>  ( .D(n18442), .E(n18285), .CK(clk), .Q(\RAM<13><1> )
         );
  EDFFX1 \RAM_reg<13><0>  ( .D(n18438), .E(n18286), .CK(clk), .Q(\RAM<13><0> )
         );
  EDFFX1 \RAM_reg<5><31>  ( .D(n18562), .E(n18300), .CK(clk), .Q(\RAM<5><31> )
         );
  EDFFX1 \RAM_reg<5><30>  ( .D(n18558), .E(n18300), .CK(clk), .Q(\RAM<5><30> )
         );
  EDFFX1 \RAM_reg<5><29>  ( .D(n18554), .E(n18300), .CK(clk), .Q(\RAM<5><29> )
         );
  EDFFX1 \RAM_reg<5><28>  ( .D(n18550), .E(n18300), .CK(clk), .Q(\RAM<5><28> )
         );
  EDFFX1 \RAM_reg<5><27>  ( .D(n18546), .E(n18300), .CK(clk), .Q(\RAM<5><27> )
         );
  EDFFX1 \RAM_reg<5><26>  ( .D(n18542), .E(n18300), .CK(clk), .Q(\RAM<5><26> )
         );
  EDFFX1 \RAM_reg<5><25>  ( .D(n18538), .E(n18300), .CK(clk), .Q(\RAM<5><25> )
         );
  EDFFX1 \RAM_reg<5><24>  ( .D(n18534), .E(n18300), .CK(clk), .Q(\RAM<5><24> )
         );
  EDFFX1 \RAM_reg<5><23>  ( .D(n18530), .E(n18300), .CK(clk), .Q(\RAM<5><23> )
         );
  EDFFX1 \RAM_reg<5><22>  ( .D(n18526), .E(n18300), .CK(clk), .Q(\RAM<5><22> )
         );
  EDFFX1 \RAM_reg<5><21>  ( .D(n18522), .E(n18300), .CK(clk), .Q(\RAM<5><21> )
         );
  EDFFX1 \RAM_reg<5><20>  ( .D(n18518), .E(n18300), .CK(clk), .Q(\RAM<5><20> )
         );
  EDFFX1 \RAM_reg<5><19>  ( .D(n18514), .E(n18301), .CK(clk), .Q(\RAM<5><19> )
         );
  EDFFX1 \RAM_reg<5><18>  ( .D(n18510), .E(n18301), .CK(clk), .Q(\RAM<5><18> )
         );
  EDFFX1 \RAM_reg<5><17>  ( .D(n18506), .E(n18301), .CK(clk), .Q(\RAM<5><17> )
         );
  EDFFX1 \RAM_reg<5><16>  ( .D(n18502), .E(n18301), .CK(clk), .Q(\RAM<5><16> )
         );
  EDFFX1 \RAM_reg<5><15>  ( .D(n18498), .E(n18301), .CK(clk), .Q(\RAM<5><15> )
         );
  EDFFX1 \RAM_reg<5><14>  ( .D(n18494), .E(n18301), .CK(clk), .Q(\RAM<5><14> )
         );
  EDFFX1 \RAM_reg<5><13>  ( .D(n18490), .E(n18301), .CK(clk), .Q(\RAM<5><13> )
         );
  EDFFX1 \RAM_reg<5><12>  ( .D(n18486), .E(n18301), .CK(clk), .Q(\RAM<5><12> )
         );
  EDFFX1 \RAM_reg<5><11>  ( .D(n18482), .E(n18301), .CK(clk), .Q(\RAM<5><11> )
         );
  EDFFX1 \RAM_reg<5><10>  ( .D(n18478), .E(n18301), .CK(clk), .Q(\RAM<5><10> )
         );
  EDFFX1 \RAM_reg<5><9>  ( .D(n18474), .E(n18301), .CK(clk), .Q(\RAM<5><9> )
         );
  EDFFX1 \RAM_reg<5><8>  ( .D(n18470), .E(n18301), .CK(clk), .Q(\RAM<5><8> )
         );
  EDFFX1 \RAM_reg<5><7>  ( .D(n18466), .E(n3570), .CK(clk), .Q(\RAM<5><7> ) );
  EDFFX1 \RAM_reg<5><6>  ( .D(n18462), .E(n3570), .CK(clk), .Q(\RAM<5><6> ) );
  EDFFX1 \RAM_reg<5><5>  ( .D(n18458), .E(n18300), .CK(clk), .Q(\RAM<5><5> )
         );
  EDFFX1 \RAM_reg<5><4>  ( .D(n18454), .E(n18301), .CK(clk), .Q(\RAM<5><4> )
         );
  EDFFX1 \RAM_reg<5><3>  ( .D(n18450), .E(n18300), .CK(clk), .Q(\RAM<5><3> )
         );
  EDFFX1 \RAM_reg<5><2>  ( .D(n18446), .E(n18301), .CK(clk), .Q(\RAM<5><2> )
         );
  EDFFX1 \RAM_reg<5><1>  ( .D(n18442), .E(n18300), .CK(clk), .Q(\RAM<5><1> )
         );
  EDFFX1 \RAM_reg<5><0>  ( .D(n18438), .E(n18301), .CK(clk), .Q(\RAM<5><0> )
         );
  EDFFX1 \RAM_reg<63><31>  ( .D(n18562), .E(n18354), .CK(clk), .Q(
        \RAM<63><31> ) );
  EDFFX1 \RAM_reg<63><30>  ( .D(n18558), .E(n18354), .CK(clk), .Q(
        \RAM<63><30> ) );
  EDFFX1 \RAM_reg<63><29>  ( .D(n18554), .E(n18354), .CK(clk), .Q(
        \RAM<63><29> ) );
  EDFFX1 \RAM_reg<63><28>  ( .D(n18550), .E(n18354), .CK(clk), .Q(
        \RAM<63><28> ) );
  EDFFX1 \RAM_reg<63><27>  ( .D(n18546), .E(n18354), .CK(clk), .Q(
        \RAM<63><27> ) );
  EDFFX1 \RAM_reg<63><26>  ( .D(n18542), .E(n18354), .CK(clk), .Q(
        \RAM<63><26> ) );
  EDFFX1 \RAM_reg<63><25>  ( .D(n18538), .E(n18354), .CK(clk), .Q(
        \RAM<63><25> ) );
  EDFFX1 \RAM_reg<63><24>  ( .D(n18534), .E(n18354), .CK(clk), .Q(
        \RAM<63><24> ) );
  EDFFX1 \RAM_reg<63><23>  ( .D(n18530), .E(n18354), .CK(clk), .Q(
        \RAM<63><23> ) );
  EDFFX1 \RAM_reg<63><22>  ( .D(n18526), .E(n18354), .CK(clk), .Q(
        \RAM<63><22> ) );
  EDFFX1 \RAM_reg<63><21>  ( .D(n18522), .E(n18354), .CK(clk), .Q(
        \RAM<63><21> ) );
  EDFFX1 \RAM_reg<63><20>  ( .D(n18518), .E(n18354), .CK(clk), .Q(
        \RAM<63><20> ) );
  EDFFX1 \RAM_reg<63><19>  ( .D(n18514), .E(n18355), .CK(clk), .Q(
        \RAM<63><19> ) );
  EDFFX1 \RAM_reg<63><18>  ( .D(n18510), .E(n18355), .CK(clk), .Q(
        \RAM<63><18> ) );
  EDFFX1 \RAM_reg<63><17>  ( .D(n18506), .E(n18355), .CK(clk), .Q(
        \RAM<63><17> ) );
  EDFFX1 \RAM_reg<63><16>  ( .D(n18502), .E(n18355), .CK(clk), .Q(
        \RAM<63><16> ) );
  EDFFX1 \RAM_reg<63><15>  ( .D(n18498), .E(n18355), .CK(clk), .Q(
        \RAM<63><15> ) );
  EDFFX1 \RAM_reg<63><14>  ( .D(n18494), .E(n18355), .CK(clk), .Q(
        \RAM<63><14> ) );
  EDFFX1 \RAM_reg<63><13>  ( .D(n18490), .E(n18355), .CK(clk), .Q(
        \RAM<63><13> ) );
  EDFFX1 \RAM_reg<63><12>  ( .D(n18486), .E(n18355), .CK(clk), .Q(
        \RAM<63><12> ) );
  EDFFX1 \RAM_reg<63><11>  ( .D(n18482), .E(n18355), .CK(clk), .Q(
        \RAM<63><11> ) );
  EDFFX1 \RAM_reg<63><10>  ( .D(n18478), .E(n18355), .CK(clk), .Q(
        \RAM<63><10> ) );
  EDFFX1 \RAM_reg<63><9>  ( .D(n18474), .E(n18355), .CK(clk), .Q(\RAM<63><9> )
         );
  EDFFX1 \RAM_reg<63><8>  ( .D(n18470), .E(n18355), .CK(clk), .Q(\RAM<63><8> )
         );
  EDFFX1 \RAM_reg<63><7>  ( .D(n18466), .E(n3546), .CK(clk), .Q(\RAM<63><7> )
         );
  EDFFX1 \RAM_reg<63><6>  ( .D(n18462), .E(n3546), .CK(clk), .Q(\RAM<63><6> )
         );
  EDFFX1 \RAM_reg<63><5>  ( .D(n18458), .E(n18354), .CK(clk), .Q(\RAM<63><5> )
         );
  EDFFX1 \RAM_reg<63><4>  ( .D(n18454), .E(n18355), .CK(clk), .Q(\RAM<63><4> )
         );
  EDFFX1 \RAM_reg<63><3>  ( .D(n18450), .E(n18354), .CK(clk), .Q(\RAM<63><3> )
         );
  EDFFX1 \RAM_reg<63><2>  ( .D(n18446), .E(n18355), .CK(clk), .Q(\RAM<63><2> )
         );
  EDFFX1 \RAM_reg<63><1>  ( .D(n18442), .E(n18354), .CK(clk), .Q(\RAM<63><1> )
         );
  EDFFX1 \RAM_reg<63><0>  ( .D(n18438), .E(n18355), .CK(clk), .Q(\RAM<63><0> )
         );
  EDFFX1 \RAM_reg<59><31>  ( .D(n18562), .E(n18360), .CK(clk), .Q(
        \RAM<59><31> ) );
  EDFFX1 \RAM_reg<59><30>  ( .D(n18558), .E(n18360), .CK(clk), .Q(
        \RAM<59><30> ) );
  EDFFX1 \RAM_reg<59><29>  ( .D(n18554), .E(n18360), .CK(clk), .Q(
        \RAM<59><29> ) );
  EDFFX1 \RAM_reg<59><28>  ( .D(n18550), .E(n18360), .CK(clk), .Q(
        \RAM<59><28> ) );
  EDFFX1 \RAM_reg<59><27>  ( .D(n18546), .E(n18360), .CK(clk), .Q(
        \RAM<59><27> ) );
  EDFFX1 \RAM_reg<59><26>  ( .D(n18542), .E(n18360), .CK(clk), .Q(
        \RAM<59><26> ) );
  EDFFX1 \RAM_reg<59><25>  ( .D(n18538), .E(n18360), .CK(clk), .Q(
        \RAM<59><25> ) );
  EDFFX1 \RAM_reg<59><24>  ( .D(n18534), .E(n18360), .CK(clk), .Q(
        \RAM<59><24> ) );
  EDFFX1 \RAM_reg<59><23>  ( .D(n18530), .E(n18360), .CK(clk), .Q(
        \RAM<59><23> ) );
  EDFFX1 \RAM_reg<59><22>  ( .D(n18526), .E(n18360), .CK(clk), .Q(
        \RAM<59><22> ) );
  EDFFX1 \RAM_reg<59><21>  ( .D(n18522), .E(n18360), .CK(clk), .Q(
        \RAM<59><21> ) );
  EDFFX1 \RAM_reg<59><20>  ( .D(n18518), .E(n18360), .CK(clk), .Q(
        \RAM<59><20> ) );
  EDFFX1 \RAM_reg<59><19>  ( .D(n18514), .E(n18361), .CK(clk), .Q(
        \RAM<59><19> ) );
  EDFFX1 \RAM_reg<59><18>  ( .D(n18510), .E(n18361), .CK(clk), .Q(
        \RAM<59><18> ) );
  EDFFX1 \RAM_reg<59><17>  ( .D(n18506), .E(n18361), .CK(clk), .Q(
        \RAM<59><17> ) );
  EDFFX1 \RAM_reg<59><16>  ( .D(n18502), .E(n18361), .CK(clk), .Q(
        \RAM<59><16> ) );
  EDFFX1 \RAM_reg<59><15>  ( .D(n18498), .E(n18361), .CK(clk), .Q(
        \RAM<59><15> ) );
  EDFFX1 \RAM_reg<59><14>  ( .D(n18494), .E(n18361), .CK(clk), .Q(
        \RAM<59><14> ) );
  EDFFX1 \RAM_reg<59><13>  ( .D(n18490), .E(n18361), .CK(clk), .Q(
        \RAM<59><13> ) );
  EDFFX1 \RAM_reg<59><12>  ( .D(n18486), .E(n18361), .CK(clk), .Q(
        \RAM<59><12> ) );
  EDFFX1 \RAM_reg<59><11>  ( .D(n18482), .E(n18361), .CK(clk), .Q(
        \RAM<59><11> ) );
  EDFFX1 \RAM_reg<59><10>  ( .D(n18478), .E(n18361), .CK(clk), .Q(
        \RAM<59><10> ) );
  EDFFX1 \RAM_reg<59><9>  ( .D(n18474), .E(n18361), .CK(clk), .Q(\RAM<59><9> )
         );
  EDFFX1 \RAM_reg<59><8>  ( .D(n18470), .E(n18361), .CK(clk), .Q(\RAM<59><8> )
         );
  EDFFX1 \RAM_reg<59><7>  ( .D(n18466), .E(n3544), .CK(clk), .Q(\RAM<59><7> )
         );
  EDFFX1 \RAM_reg<59><6>  ( .D(n18462), .E(n3544), .CK(clk), .Q(\RAM<59><6> )
         );
  EDFFX1 \RAM_reg<59><5>  ( .D(n18458), .E(n18360), .CK(clk), .Q(\RAM<59><5> )
         );
  EDFFX1 \RAM_reg<59><4>  ( .D(n18454), .E(n18361), .CK(clk), .Q(\RAM<59><4> )
         );
  EDFFX1 \RAM_reg<59><3>  ( .D(n18450), .E(n18360), .CK(clk), .Q(\RAM<59><3> )
         );
  EDFFX1 \RAM_reg<59><2>  ( .D(n18446), .E(n18361), .CK(clk), .Q(\RAM<59><2> )
         );
  EDFFX1 \RAM_reg<59><1>  ( .D(n18442), .E(n18360), .CK(clk), .Q(\RAM<59><1> )
         );
  EDFFX1 \RAM_reg<59><0>  ( .D(n18438), .E(n18361), .CK(clk), .Q(\RAM<59><0> )
         );
  EDFFX1 \RAM_reg<55><31>  ( .D(n18562), .E(n18351), .CK(clk), .Q(
        \RAM<55><31> ) );
  EDFFX1 \RAM_reg<55><30>  ( .D(n18558), .E(n18351), .CK(clk), .Q(
        \RAM<55><30> ) );
  EDFFX1 \RAM_reg<55><29>  ( .D(n18554), .E(n18351), .CK(clk), .Q(
        \RAM<55><29> ) );
  EDFFX1 \RAM_reg<55><28>  ( .D(n18550), .E(n18351), .CK(clk), .Q(
        \RAM<55><28> ) );
  EDFFX1 \RAM_reg<55><27>  ( .D(n18546), .E(n18351), .CK(clk), .Q(
        \RAM<55><27> ) );
  EDFFX1 \RAM_reg<55><26>  ( .D(n18542), .E(n18351), .CK(clk), .Q(
        \RAM<55><26> ) );
  EDFFX1 \RAM_reg<55><25>  ( .D(n18538), .E(n18351), .CK(clk), .Q(
        \RAM<55><25> ) );
  EDFFX1 \RAM_reg<55><24>  ( .D(n18534), .E(n18351), .CK(clk), .Q(
        \RAM<55><24> ) );
  EDFFX1 \RAM_reg<55><23>  ( .D(n18530), .E(n18351), .CK(clk), .Q(
        \RAM<55><23> ) );
  EDFFX1 \RAM_reg<55><22>  ( .D(n18526), .E(n18351), .CK(clk), .Q(
        \RAM<55><22> ) );
  EDFFX1 \RAM_reg<55><21>  ( .D(n18522), .E(n18351), .CK(clk), .Q(
        \RAM<55><21> ) );
  EDFFX1 \RAM_reg<55><20>  ( .D(n18518), .E(n18351), .CK(clk), .Q(
        \RAM<55><20> ) );
  EDFFX1 \RAM_reg<55><19>  ( .D(n18514), .E(n18352), .CK(clk), .Q(
        \RAM<55><19> ) );
  EDFFX1 \RAM_reg<55><18>  ( .D(n18510), .E(n18352), .CK(clk), .Q(
        \RAM<55><18> ) );
  EDFFX1 \RAM_reg<55><17>  ( .D(n18506), .E(n18352), .CK(clk), .Q(
        \RAM<55><17> ) );
  EDFFX1 \RAM_reg<55><16>  ( .D(n18502), .E(n18352), .CK(clk), .Q(
        \RAM<55><16> ) );
  EDFFX1 \RAM_reg<55><15>  ( .D(n18498), .E(n18352), .CK(clk), .Q(
        \RAM<55><15> ) );
  EDFFX1 \RAM_reg<55><14>  ( .D(n18494), .E(n18352), .CK(clk), .Q(
        \RAM<55><14> ) );
  EDFFX1 \RAM_reg<55><13>  ( .D(n18490), .E(n18352), .CK(clk), .Q(
        \RAM<55><13> ) );
  EDFFX1 \RAM_reg<55><12>  ( .D(n18486), .E(n18352), .CK(clk), .Q(
        \RAM<55><12> ) );
  EDFFX1 \RAM_reg<55><11>  ( .D(n18482), .E(n18352), .CK(clk), .Q(
        \RAM<55><11> ) );
  EDFFX1 \RAM_reg<55><10>  ( .D(n18478), .E(n18352), .CK(clk), .Q(
        \RAM<55><10> ) );
  EDFFX1 \RAM_reg<55><9>  ( .D(n18474), .E(n18352), .CK(clk), .Q(\RAM<55><9> )
         );
  EDFFX1 \RAM_reg<55><8>  ( .D(n18470), .E(n18352), .CK(clk), .Q(\RAM<55><8> )
         );
  EDFFX1 \RAM_reg<55><7>  ( .D(n18466), .E(n3548), .CK(clk), .Q(\RAM<55><7> )
         );
  EDFFX1 \RAM_reg<55><6>  ( .D(n18462), .E(n3548), .CK(clk), .Q(\RAM<55><6> )
         );
  EDFFX1 \RAM_reg<55><5>  ( .D(n18458), .E(n18351), .CK(clk), .Q(\RAM<55><5> )
         );
  EDFFX1 \RAM_reg<55><4>  ( .D(n18454), .E(n18352), .CK(clk), .Q(\RAM<55><4> )
         );
  EDFFX1 \RAM_reg<55><3>  ( .D(n18450), .E(n18351), .CK(clk), .Q(\RAM<55><3> )
         );
  EDFFX1 \RAM_reg<55><2>  ( .D(n18446), .E(n18352), .CK(clk), .Q(\RAM<55><2> )
         );
  EDFFX1 \RAM_reg<55><1>  ( .D(n18442), .E(n18351), .CK(clk), .Q(\RAM<55><1> )
         );
  EDFFX1 \RAM_reg<55><0>  ( .D(n18438), .E(n18352), .CK(clk), .Q(\RAM<55><0> )
         );
  EDFFX1 \RAM_reg<51><31>  ( .D(n18562), .E(n18321), .CK(clk), .Q(
        \RAM<51><31> ) );
  EDFFX1 \RAM_reg<51><30>  ( .D(n18558), .E(n18321), .CK(clk), .Q(
        \RAM<51><30> ) );
  EDFFX1 \RAM_reg<51><29>  ( .D(n18554), .E(n18321), .CK(clk), .Q(
        \RAM<51><29> ) );
  EDFFX1 \RAM_reg<51><28>  ( .D(n18550), .E(n18321), .CK(clk), .Q(
        \RAM<51><28> ) );
  EDFFX1 \RAM_reg<51><27>  ( .D(n18546), .E(n18321), .CK(clk), .Q(
        \RAM<51><27> ) );
  EDFFX1 \RAM_reg<51><26>  ( .D(n18542), .E(n18321), .CK(clk), .Q(
        \RAM<51><26> ) );
  EDFFX1 \RAM_reg<51><25>  ( .D(n18538), .E(n18321), .CK(clk), .Q(
        \RAM<51><25> ) );
  EDFFX1 \RAM_reg<51><24>  ( .D(n18534), .E(n18321), .CK(clk), .Q(
        \RAM<51><24> ) );
  EDFFX1 \RAM_reg<51><23>  ( .D(n18530), .E(n18321), .CK(clk), .Q(
        \RAM<51><23> ) );
  EDFFX1 \RAM_reg<51><22>  ( .D(n18526), .E(n18321), .CK(clk), .Q(
        \RAM<51><22> ) );
  EDFFX1 \RAM_reg<51><21>  ( .D(n18522), .E(n18321), .CK(clk), .Q(
        \RAM<51><21> ) );
  EDFFX1 \RAM_reg<51><20>  ( .D(n18518), .E(n18321), .CK(clk), .Q(
        \RAM<51><20> ) );
  EDFFX1 \RAM_reg<51><19>  ( .D(n18514), .E(n18322), .CK(clk), .Q(
        \RAM<51><19> ) );
  EDFFX1 \RAM_reg<51><18>  ( .D(n18510), .E(n18322), .CK(clk), .Q(
        \RAM<51><18> ) );
  EDFFX1 \RAM_reg<51><17>  ( .D(n18506), .E(n18322), .CK(clk), .Q(
        \RAM<51><17> ) );
  EDFFX1 \RAM_reg<51><16>  ( .D(n18502), .E(n18322), .CK(clk), .Q(
        \RAM<51><16> ) );
  EDFFX1 \RAM_reg<51><15>  ( .D(n18498), .E(n18322), .CK(clk), .Q(
        \RAM<51><15> ) );
  EDFFX1 \RAM_reg<51><14>  ( .D(n18494), .E(n18322), .CK(clk), .Q(
        \RAM<51><14> ) );
  EDFFX1 \RAM_reg<51><13>  ( .D(n18490), .E(n18322), .CK(clk), .Q(
        \RAM<51><13> ) );
  EDFFX1 \RAM_reg<51><12>  ( .D(n18486), .E(n18322), .CK(clk), .Q(
        \RAM<51><12> ) );
  EDFFX1 \RAM_reg<51><11>  ( .D(n18482), .E(n18322), .CK(clk), .Q(
        \RAM<51><11> ) );
  EDFFX1 \RAM_reg<51><10>  ( .D(n18478), .E(n18322), .CK(clk), .Q(
        \RAM<51><10> ) );
  EDFFX1 \RAM_reg<51><9>  ( .D(n18474), .E(n18322), .CK(clk), .Q(\RAM<51><9> )
         );
  EDFFX1 \RAM_reg<51><8>  ( .D(n18470), .E(n18322), .CK(clk), .Q(\RAM<51><8> )
         );
  EDFFX1 \RAM_reg<51><7>  ( .D(n18466), .E(n3558), .CK(clk), .Q(\RAM<51><7> )
         );
  EDFFX1 \RAM_reg<51><6>  ( .D(n18462), .E(n3558), .CK(clk), .Q(\RAM<51><6> )
         );
  EDFFX1 \RAM_reg<51><5>  ( .D(n18458), .E(n18321), .CK(clk), .Q(\RAM<51><5> )
         );
  EDFFX1 \RAM_reg<51><4>  ( .D(n18454), .E(n18322), .CK(clk), .Q(\RAM<51><4> )
         );
  EDFFX1 \RAM_reg<51><3>  ( .D(n18450), .E(n18321), .CK(clk), .Q(\RAM<51><3> )
         );
  EDFFX1 \RAM_reg<51><2>  ( .D(n18446), .E(n18322), .CK(clk), .Q(\RAM<51><2> )
         );
  EDFFX1 \RAM_reg<51><1>  ( .D(n18442), .E(n18321), .CK(clk), .Q(\RAM<51><1> )
         );
  EDFFX1 \RAM_reg<51><0>  ( .D(n18438), .E(n18322), .CK(clk), .Q(\RAM<51><0> )
         );
  EDFFX1 \RAM_reg<47><31>  ( .D(n18563), .E(n18405), .CK(clk), .Q(
        \RAM<47><31> ) );
  EDFFX1 \RAM_reg<47><30>  ( .D(n18559), .E(n18405), .CK(clk), .Q(
        \RAM<47><30> ) );
  EDFFX1 \RAM_reg<47><29>  ( .D(n18555), .E(n18405), .CK(clk), .Q(
        \RAM<47><29> ) );
  EDFFX1 \RAM_reg<47><28>  ( .D(n18551), .E(n18405), .CK(clk), .Q(
        \RAM<47><28> ) );
  EDFFX1 \RAM_reg<47><27>  ( .D(n18547), .E(n18405), .CK(clk), .Q(
        \RAM<47><27> ) );
  EDFFX1 \RAM_reg<47><26>  ( .D(n18543), .E(n18405), .CK(clk), .Q(
        \RAM<47><26> ) );
  EDFFX1 \RAM_reg<47><25>  ( .D(n18539), .E(n18405), .CK(clk), .Q(
        \RAM<47><25> ) );
  EDFFX1 \RAM_reg<47><24>  ( .D(n18535), .E(n18405), .CK(clk), .Q(
        \RAM<47><24> ) );
  EDFFX1 \RAM_reg<47><23>  ( .D(n18531), .E(n18405), .CK(clk), .Q(
        \RAM<47><23> ) );
  EDFFX1 \RAM_reg<47><22>  ( .D(n18527), .E(n18405), .CK(clk), .Q(
        \RAM<47><22> ) );
  EDFFX1 \RAM_reg<47><21>  ( .D(n18523), .E(n18405), .CK(clk), .Q(
        \RAM<47><21> ) );
  EDFFX1 \RAM_reg<47><20>  ( .D(n18519), .E(n18405), .CK(clk), .Q(
        \RAM<47><20> ) );
  EDFFX1 \RAM_reg<47><19>  ( .D(n18515), .E(n18406), .CK(clk), .Q(
        \RAM<47><19> ) );
  EDFFX1 \RAM_reg<47><18>  ( .D(n18511), .E(n18406), .CK(clk), .Q(
        \RAM<47><18> ) );
  EDFFX1 \RAM_reg<47><17>  ( .D(n18507), .E(n18406), .CK(clk), .Q(
        \RAM<47><17> ) );
  EDFFX1 \RAM_reg<47><16>  ( .D(n18503), .E(n18406), .CK(clk), .Q(
        \RAM<47><16> ) );
  EDFFX1 \RAM_reg<47><15>  ( .D(n18499), .E(n18406), .CK(clk), .Q(
        \RAM<47><15> ) );
  EDFFX1 \RAM_reg<47><14>  ( .D(n18495), .E(n18406), .CK(clk), .Q(
        \RAM<47><14> ) );
  EDFFX1 \RAM_reg<47><13>  ( .D(n18491), .E(n18406), .CK(clk), .Q(
        \RAM<47><13> ) );
  EDFFX1 \RAM_reg<47><12>  ( .D(n18487), .E(n18406), .CK(clk), .Q(
        \RAM<47><12> ) );
  EDFFX1 \RAM_reg<47><11>  ( .D(n18483), .E(n18406), .CK(clk), .Q(
        \RAM<47><11> ) );
  EDFFX1 \RAM_reg<47><10>  ( .D(n18479), .E(n18406), .CK(clk), .Q(
        \RAM<47><10> ) );
  EDFFX1 \RAM_reg<47><9>  ( .D(n18475), .E(n18406), .CK(clk), .Q(\RAM<47><9> )
         );
  EDFFX1 \RAM_reg<47><8>  ( .D(n18471), .E(n18406), .CK(clk), .Q(\RAM<47><8> )
         );
  EDFFX1 \RAM_reg<47><7>  ( .D(n18467), .E(n3528), .CK(clk), .Q(\RAM<47><7> )
         );
  EDFFX1 \RAM_reg<47><6>  ( .D(n18463), .E(n3528), .CK(clk), .Q(\RAM<47><6> )
         );
  EDFFX1 \RAM_reg<47><5>  ( .D(n18459), .E(n18405), .CK(clk), .Q(\RAM<47><5> )
         );
  EDFFX1 \RAM_reg<47><4>  ( .D(n18455), .E(n18406), .CK(clk), .Q(\RAM<47><4> )
         );
  EDFFX1 \RAM_reg<47><3>  ( .D(n18451), .E(n18405), .CK(clk), .Q(\RAM<47><3> )
         );
  EDFFX1 \RAM_reg<47><2>  ( .D(n18447), .E(n18406), .CK(clk), .Q(\RAM<47><2> )
         );
  EDFFX1 \RAM_reg<47><1>  ( .D(n18443), .E(n18405), .CK(clk), .Q(\RAM<47><1> )
         );
  EDFFX1 \RAM_reg<47><0>  ( .D(n18439), .E(n18406), .CK(clk), .Q(\RAM<47><0> )
         );
  EDFFX1 \RAM_reg<43><31>  ( .D(n18563), .E(n18402), .CK(clk), .Q(
        \RAM<43><31> ) );
  EDFFX1 \RAM_reg<43><30>  ( .D(n18559), .E(n18402), .CK(clk), .Q(
        \RAM<43><30> ) );
  EDFFX1 \RAM_reg<43><29>  ( .D(n18555), .E(n18402), .CK(clk), .Q(
        \RAM<43><29> ) );
  EDFFX1 \RAM_reg<43><28>  ( .D(n18551), .E(n18402), .CK(clk), .Q(
        \RAM<43><28> ) );
  EDFFX1 \RAM_reg<43><27>  ( .D(n18547), .E(n18402), .CK(clk), .Q(
        \RAM<43><27> ) );
  EDFFX1 \RAM_reg<43><26>  ( .D(n18543), .E(n18402), .CK(clk), .Q(
        \RAM<43><26> ) );
  EDFFX1 \RAM_reg<43><25>  ( .D(n18539), .E(n18402), .CK(clk), .Q(
        \RAM<43><25> ) );
  EDFFX1 \RAM_reg<43><24>  ( .D(n18535), .E(n18402), .CK(clk), .Q(
        \RAM<43><24> ) );
  EDFFX1 \RAM_reg<43><23>  ( .D(n18531), .E(n18402), .CK(clk), .Q(
        \RAM<43><23> ) );
  EDFFX1 \RAM_reg<43><22>  ( .D(n18527), .E(n18402), .CK(clk), .Q(
        \RAM<43><22> ) );
  EDFFX1 \RAM_reg<43><21>  ( .D(n18523), .E(n18402), .CK(clk), .Q(
        \RAM<43><21> ) );
  EDFFX1 \RAM_reg<43><20>  ( .D(n18519), .E(n18402), .CK(clk), .Q(
        \RAM<43><20> ) );
  EDFFX1 \RAM_reg<43><19>  ( .D(n18515), .E(n18403), .CK(clk), .Q(
        \RAM<43><19> ) );
  EDFFX1 \RAM_reg<43><18>  ( .D(n18511), .E(n18403), .CK(clk), .Q(
        \RAM<43><18> ) );
  EDFFX1 \RAM_reg<43><17>  ( .D(n18507), .E(n18403), .CK(clk), .Q(
        \RAM<43><17> ) );
  EDFFX1 \RAM_reg<43><16>  ( .D(n18503), .E(n18403), .CK(clk), .Q(
        \RAM<43><16> ) );
  EDFFX1 \RAM_reg<43><15>  ( .D(n18499), .E(n18403), .CK(clk), .Q(
        \RAM<43><15> ) );
  EDFFX1 \RAM_reg<43><14>  ( .D(n18495), .E(n18403), .CK(clk), .Q(
        \RAM<43><14> ) );
  EDFFX1 \RAM_reg<43><13>  ( .D(n18491), .E(n18403), .CK(clk), .Q(
        \RAM<43><13> ) );
  EDFFX1 \RAM_reg<43><12>  ( .D(n18487), .E(n18403), .CK(clk), .Q(
        \RAM<43><12> ) );
  EDFFX1 \RAM_reg<43><11>  ( .D(n18483), .E(n18403), .CK(clk), .Q(
        \RAM<43><11> ) );
  EDFFX1 \RAM_reg<43><10>  ( .D(n18479), .E(n18403), .CK(clk), .Q(
        \RAM<43><10> ) );
  EDFFX1 \RAM_reg<43><9>  ( .D(n18475), .E(n18403), .CK(clk), .Q(\RAM<43><9> )
         );
  EDFFX1 \RAM_reg<43><8>  ( .D(n18471), .E(n18403), .CK(clk), .Q(\RAM<43><8> )
         );
  EDFFX1 \RAM_reg<43><7>  ( .D(n18467), .E(n3529), .CK(clk), .Q(\RAM<43><7> )
         );
  EDFFX1 \RAM_reg<43><6>  ( .D(n18463), .E(n3529), .CK(clk), .Q(\RAM<43><6> )
         );
  EDFFX1 \RAM_reg<43><5>  ( .D(n18459), .E(n18402), .CK(clk), .Q(\RAM<43><5> )
         );
  EDFFX1 \RAM_reg<43><4>  ( .D(n18455), .E(n18403), .CK(clk), .Q(\RAM<43><4> )
         );
  EDFFX1 \RAM_reg<43><3>  ( .D(n18451), .E(n18402), .CK(clk), .Q(\RAM<43><3> )
         );
  EDFFX1 \RAM_reg<43><2>  ( .D(n18447), .E(n18403), .CK(clk), .Q(\RAM<43><2> )
         );
  EDFFX1 \RAM_reg<43><1>  ( .D(n18443), .E(n18402), .CK(clk), .Q(\RAM<43><1> )
         );
  EDFFX1 \RAM_reg<43><0>  ( .D(n18439), .E(n18403), .CK(clk), .Q(\RAM<43><0> )
         );
  EDFFX1 \RAM_reg<39><31>  ( .D(n18563), .E(n18408), .CK(clk), .Q(
        \RAM<39><31> ) );
  EDFFX1 \RAM_reg<39><30>  ( .D(n18559), .E(n18408), .CK(clk), .Q(
        \RAM<39><30> ) );
  EDFFX1 \RAM_reg<39><29>  ( .D(n18555), .E(n18408), .CK(clk), .Q(
        \RAM<39><29> ) );
  EDFFX1 \RAM_reg<39><28>  ( .D(n18551), .E(n18408), .CK(clk), .Q(
        \RAM<39><28> ) );
  EDFFX1 \RAM_reg<39><27>  ( .D(n18547), .E(n18408), .CK(clk), .Q(
        \RAM<39><27> ) );
  EDFFX1 \RAM_reg<39><26>  ( .D(n18543), .E(n18408), .CK(clk), .Q(
        \RAM<39><26> ) );
  EDFFX1 \RAM_reg<39><25>  ( .D(n18539), .E(n18408), .CK(clk), .Q(
        \RAM<39><25> ) );
  EDFFX1 \RAM_reg<39><24>  ( .D(n18535), .E(n18408), .CK(clk), .Q(
        \RAM<39><24> ) );
  EDFFX1 \RAM_reg<39><23>  ( .D(n18531), .E(n18408), .CK(clk), .Q(
        \RAM<39><23> ) );
  EDFFX1 \RAM_reg<39><22>  ( .D(n18527), .E(n18408), .CK(clk), .Q(
        \RAM<39><22> ) );
  EDFFX1 \RAM_reg<39><21>  ( .D(n18523), .E(n18408), .CK(clk), .Q(
        \RAM<39><21> ) );
  EDFFX1 \RAM_reg<39><20>  ( .D(n18519), .E(n18408), .CK(clk), .Q(
        \RAM<39><20> ) );
  EDFFX1 \RAM_reg<39><19>  ( .D(n18515), .E(n18409), .CK(clk), .Q(
        \RAM<39><19> ) );
  EDFFX1 \RAM_reg<39><18>  ( .D(n18511), .E(n18409), .CK(clk), .Q(
        \RAM<39><18> ) );
  EDFFX1 \RAM_reg<39><17>  ( .D(n18507), .E(n18409), .CK(clk), .Q(
        \RAM<39><17> ) );
  EDFFX1 \RAM_reg<39><16>  ( .D(n18503), .E(n18409), .CK(clk), .Q(
        \RAM<39><16> ) );
  EDFFX1 \RAM_reg<39><15>  ( .D(n18499), .E(n18409), .CK(clk), .Q(
        \RAM<39><15> ) );
  EDFFX1 \RAM_reg<39><14>  ( .D(n18495), .E(n18409), .CK(clk), .Q(
        \RAM<39><14> ) );
  EDFFX1 \RAM_reg<39><13>  ( .D(n18491), .E(n18409), .CK(clk), .Q(
        \RAM<39><13> ) );
  EDFFX1 \RAM_reg<39><12>  ( .D(n18487), .E(n18409), .CK(clk), .Q(
        \RAM<39><12> ) );
  EDFFX1 \RAM_reg<39><11>  ( .D(n18483), .E(n18409), .CK(clk), .Q(
        \RAM<39><11> ) );
  EDFFX1 \RAM_reg<39><10>  ( .D(n18479), .E(n18409), .CK(clk), .Q(
        \RAM<39><10> ) );
  EDFFX1 \RAM_reg<39><9>  ( .D(n18475), .E(n18409), .CK(clk), .Q(\RAM<39><9> )
         );
  EDFFX1 \RAM_reg<39><8>  ( .D(n18471), .E(n18409), .CK(clk), .Q(\RAM<39><8> )
         );
  EDFFX1 \RAM_reg<39><7>  ( .D(n18467), .E(n3527), .CK(clk), .Q(\RAM<39><7> )
         );
  EDFFX1 \RAM_reg<39><6>  ( .D(n18463), .E(n3527), .CK(clk), .Q(\RAM<39><6> )
         );
  EDFFX1 \RAM_reg<39><5>  ( .D(n18459), .E(n18408), .CK(clk), .Q(\RAM<39><5> )
         );
  EDFFX1 \RAM_reg<39><4>  ( .D(n18455), .E(n18409), .CK(clk), .Q(\RAM<39><4> )
         );
  EDFFX1 \RAM_reg<39><3>  ( .D(n18451), .E(n18408), .CK(clk), .Q(\RAM<39><3> )
         );
  EDFFX1 \RAM_reg<39><2>  ( .D(n18447), .E(n18409), .CK(clk), .Q(\RAM<39><2> )
         );
  EDFFX1 \RAM_reg<39><1>  ( .D(n18443), .E(n18408), .CK(clk), .Q(\RAM<39><1> )
         );
  EDFFX1 \RAM_reg<39><0>  ( .D(n18439), .E(n18409), .CK(clk), .Q(\RAM<39><0> )
         );
  EDFFX1 \RAM_reg<35><31>  ( .D(n18563), .E(n18399), .CK(clk), .Q(
        \RAM<35><31> ) );
  EDFFX1 \RAM_reg<35><30>  ( .D(n18559), .E(n18399), .CK(clk), .Q(
        \RAM<35><30> ) );
  EDFFX1 \RAM_reg<35><29>  ( .D(n18555), .E(n18399), .CK(clk), .Q(
        \RAM<35><29> ) );
  EDFFX1 \RAM_reg<35><28>  ( .D(n18551), .E(n18399), .CK(clk), .Q(
        \RAM<35><28> ) );
  EDFFX1 \RAM_reg<35><27>  ( .D(n18547), .E(n18399), .CK(clk), .Q(
        \RAM<35><27> ) );
  EDFFX1 \RAM_reg<35><26>  ( .D(n18543), .E(n18399), .CK(clk), .Q(
        \RAM<35><26> ) );
  EDFFX1 \RAM_reg<35><25>  ( .D(n18539), .E(n18399), .CK(clk), .Q(
        \RAM<35><25> ) );
  EDFFX1 \RAM_reg<35><24>  ( .D(n18535), .E(n18399), .CK(clk), .Q(
        \RAM<35><24> ) );
  EDFFX1 \RAM_reg<35><23>  ( .D(n18531), .E(n18399), .CK(clk), .Q(
        \RAM<35><23> ) );
  EDFFX1 \RAM_reg<35><22>  ( .D(n18527), .E(n18399), .CK(clk), .Q(
        \RAM<35><22> ) );
  EDFFX1 \RAM_reg<35><21>  ( .D(n18523), .E(n18399), .CK(clk), .Q(
        \RAM<35><21> ) );
  EDFFX1 \RAM_reg<35><20>  ( .D(n18519), .E(n18399), .CK(clk), .Q(
        \RAM<35><20> ) );
  EDFFX1 \RAM_reg<35><19>  ( .D(n18515), .E(n18400), .CK(clk), .Q(
        \RAM<35><19> ) );
  EDFFX1 \RAM_reg<35><18>  ( .D(n18511), .E(n18400), .CK(clk), .Q(
        \RAM<35><18> ) );
  EDFFX1 \RAM_reg<35><17>  ( .D(n18507), .E(n18400), .CK(clk), .Q(
        \RAM<35><17> ) );
  EDFFX1 \RAM_reg<35><16>  ( .D(n18503), .E(n18400), .CK(clk), .Q(
        \RAM<35><16> ) );
  EDFFX1 \RAM_reg<35><15>  ( .D(n18499), .E(n18400), .CK(clk), .Q(
        \RAM<35><15> ) );
  EDFFX1 \RAM_reg<35><14>  ( .D(n18495), .E(n18400), .CK(clk), .Q(
        \RAM<35><14> ) );
  EDFFX1 \RAM_reg<35><13>  ( .D(n18491), .E(n18400), .CK(clk), .Q(
        \RAM<35><13> ) );
  EDFFX1 \RAM_reg<35><12>  ( .D(n18487), .E(n18400), .CK(clk), .Q(
        \RAM<35><12> ) );
  EDFFX1 \RAM_reg<35><11>  ( .D(n18483), .E(n18400), .CK(clk), .Q(
        \RAM<35><11> ) );
  EDFFX1 \RAM_reg<35><10>  ( .D(n18479), .E(n18400), .CK(clk), .Q(
        \RAM<35><10> ) );
  EDFFX1 \RAM_reg<35><9>  ( .D(n18475), .E(n18400), .CK(clk), .Q(\RAM<35><9> )
         );
  EDFFX1 \RAM_reg<35><8>  ( .D(n18471), .E(n18400), .CK(clk), .Q(\RAM<35><8> )
         );
  EDFFX1 \RAM_reg<35><7>  ( .D(n18467), .E(n3530), .CK(clk), .Q(\RAM<35><7> )
         );
  EDFFX1 \RAM_reg<35><6>  ( .D(n18463), .E(n3530), .CK(clk), .Q(\RAM<35><6> )
         );
  EDFFX1 \RAM_reg<35><5>  ( .D(n18459), .E(n18399), .CK(clk), .Q(\RAM<35><5> )
         );
  EDFFX1 \RAM_reg<35><4>  ( .D(n18455), .E(n18400), .CK(clk), .Q(\RAM<35><4> )
         );
  EDFFX1 \RAM_reg<35><3>  ( .D(n18451), .E(n18399), .CK(clk), .Q(\RAM<35><3> )
         );
  EDFFX1 \RAM_reg<35><2>  ( .D(n18447), .E(n18400), .CK(clk), .Q(\RAM<35><2> )
         );
  EDFFX1 \RAM_reg<35><1>  ( .D(n18443), .E(n18399), .CK(clk), .Q(\RAM<35><1> )
         );
  EDFFX1 \RAM_reg<35><0>  ( .D(n18439), .E(n18400), .CK(clk), .Q(\RAM<35><0> )
         );
  EDFFX1 \RAM_reg<31><31>  ( .D(n18563), .E(n18378), .CK(clk), .Q(
        \RAM<31><31> ) );
  EDFFX1 \RAM_reg<31><30>  ( .D(n18559), .E(n18378), .CK(clk), .Q(
        \RAM<31><30> ) );
  EDFFX1 \RAM_reg<31><29>  ( .D(n18555), .E(n18378), .CK(clk), .Q(
        \RAM<31><29> ) );
  EDFFX1 \RAM_reg<31><28>  ( .D(n18551), .E(n18378), .CK(clk), .Q(
        \RAM<31><28> ) );
  EDFFX1 \RAM_reg<31><27>  ( .D(n18547), .E(n18378), .CK(clk), .Q(
        \RAM<31><27> ) );
  EDFFX1 \RAM_reg<31><26>  ( .D(n18543), .E(n18378), .CK(clk), .Q(
        \RAM<31><26> ) );
  EDFFX1 \RAM_reg<31><25>  ( .D(n18539), .E(n18378), .CK(clk), .Q(
        \RAM<31><25> ) );
  EDFFX1 \RAM_reg<31><24>  ( .D(n18535), .E(n18378), .CK(clk), .Q(
        \RAM<31><24> ) );
  EDFFX1 \RAM_reg<31><23>  ( .D(n18531), .E(n18378), .CK(clk), .Q(
        \RAM<31><23> ) );
  EDFFX1 \RAM_reg<31><22>  ( .D(n18527), .E(n18378), .CK(clk), .Q(
        \RAM<31><22> ) );
  EDFFX1 \RAM_reg<31><21>  ( .D(n18523), .E(n18378), .CK(clk), .Q(
        \RAM<31><21> ) );
  EDFFX1 \RAM_reg<31><20>  ( .D(n18519), .E(n18378), .CK(clk), .Q(
        \RAM<31><20> ) );
  EDFFX1 \RAM_reg<31><19>  ( .D(n18515), .E(n18379), .CK(clk), .Q(
        \RAM<31><19> ) );
  EDFFX1 \RAM_reg<31><18>  ( .D(n18511), .E(n18379), .CK(clk), .Q(
        \RAM<31><18> ) );
  EDFFX1 \RAM_reg<31><17>  ( .D(n18507), .E(n18379), .CK(clk), .Q(
        \RAM<31><17> ) );
  EDFFX1 \RAM_reg<31><16>  ( .D(n18503), .E(n18379), .CK(clk), .Q(
        \RAM<31><16> ) );
  EDFFX1 \RAM_reg<31><15>  ( .D(n18499), .E(n18379), .CK(clk), .Q(
        \RAM<31><15> ) );
  EDFFX1 \RAM_reg<31><14>  ( .D(n18495), .E(n18379), .CK(clk), .Q(
        \RAM<31><14> ) );
  EDFFX1 \RAM_reg<31><13>  ( .D(n18491), .E(n18379), .CK(clk), .Q(
        \RAM<31><13> ) );
  EDFFX1 \RAM_reg<31><12>  ( .D(n18487), .E(n18379), .CK(clk), .Q(
        \RAM<31><12> ) );
  EDFFX1 \RAM_reg<31><11>  ( .D(n18483), .E(n18379), .CK(clk), .Q(
        \RAM<31><11> ) );
  EDFFX1 \RAM_reg<31><10>  ( .D(n18479), .E(n18379), .CK(clk), .Q(
        \RAM<31><10> ) );
  EDFFX1 \RAM_reg<31><9>  ( .D(n18475), .E(n18379), .CK(clk), .Q(\RAM<31><9> )
         );
  EDFFX1 \RAM_reg<31><8>  ( .D(n18471), .E(n18379), .CK(clk), .Q(\RAM<31><8> )
         );
  EDFFX1 \RAM_reg<31><7>  ( .D(n18467), .E(n3538), .CK(clk), .Q(\RAM<31><7> )
         );
  EDFFX1 \RAM_reg<31><6>  ( .D(n18463), .E(n3538), .CK(clk), .Q(\RAM<31><6> )
         );
  EDFFX1 \RAM_reg<31><5>  ( .D(n18459), .E(n18378), .CK(clk), .Q(\RAM<31><5> )
         );
  EDFFX1 \RAM_reg<31><4>  ( .D(n18455), .E(n18379), .CK(clk), .Q(\RAM<31><4> )
         );
  EDFFX1 \RAM_reg<31><3>  ( .D(n18451), .E(n18378), .CK(clk), .Q(\RAM<31><3> )
         );
  EDFFX1 \RAM_reg<31><2>  ( .D(n18447), .E(n18379), .CK(clk), .Q(\RAM<31><2> )
         );
  EDFFX1 \RAM_reg<31><1>  ( .D(n18443), .E(n18378), .CK(clk), .Q(\RAM<31><1> )
         );
  EDFFX1 \RAM_reg<31><0>  ( .D(n18439), .E(n18379), .CK(clk), .Q(\RAM<31><0> )
         );
  EDFFX1 \RAM_reg<27><31>  ( .D(n18563), .E(n18420), .CK(clk), .Q(
        \RAM<27><31> ) );
  EDFFX1 \RAM_reg<27><30>  ( .D(n18559), .E(n18420), .CK(clk), .Q(
        \RAM<27><30> ) );
  EDFFX1 \RAM_reg<27><29>  ( .D(n18555), .E(n18420), .CK(clk), .Q(
        \RAM<27><29> ) );
  EDFFX1 \RAM_reg<27><28>  ( .D(n18551), .E(n18420), .CK(clk), .Q(
        \RAM<27><28> ) );
  EDFFX1 \RAM_reg<27><27>  ( .D(n18547), .E(n18420), .CK(clk), .Q(
        \RAM<27><27> ) );
  EDFFX1 \RAM_reg<27><26>  ( .D(n18543), .E(n18420), .CK(clk), .Q(
        \RAM<27><26> ) );
  EDFFX1 \RAM_reg<27><25>  ( .D(n18539), .E(n18420), .CK(clk), .Q(
        \RAM<27><25> ) );
  EDFFX1 \RAM_reg<27><24>  ( .D(n18535), .E(n18420), .CK(clk), .Q(
        \RAM<27><24> ) );
  EDFFX1 \RAM_reg<27><23>  ( .D(n18531), .E(n18420), .CK(clk), .Q(
        \RAM<27><23> ) );
  EDFFX1 \RAM_reg<27><22>  ( .D(n18527), .E(n18420), .CK(clk), .Q(
        \RAM<27><22> ) );
  EDFFX1 \RAM_reg<27><21>  ( .D(n18523), .E(n18420), .CK(clk), .Q(
        \RAM<27><21> ) );
  EDFFX1 \RAM_reg<27><20>  ( .D(n18519), .E(n18420), .CK(clk), .Q(
        \RAM<27><20> ) );
  EDFFX1 \RAM_reg<27><19>  ( .D(n18515), .E(n18421), .CK(clk), .Q(
        \RAM<27><19> ) );
  EDFFX1 \RAM_reg<27><18>  ( .D(n18511), .E(n18421), .CK(clk), .Q(
        \RAM<27><18> ) );
  EDFFX1 \RAM_reg<27><17>  ( .D(n18507), .E(n18421), .CK(clk), .Q(
        \RAM<27><17> ) );
  EDFFX1 \RAM_reg<27><16>  ( .D(n18503), .E(n18421), .CK(clk), .Q(
        \RAM<27><16> ) );
  EDFFX1 \RAM_reg<27><15>  ( .D(n18499), .E(n18421), .CK(clk), .Q(
        \RAM<27><15> ) );
  EDFFX1 \RAM_reg<27><14>  ( .D(n18495), .E(n18421), .CK(clk), .Q(
        \RAM<27><14> ) );
  EDFFX1 \RAM_reg<27><13>  ( .D(n18491), .E(n18421), .CK(clk), .Q(
        \RAM<27><13> ) );
  EDFFX1 \RAM_reg<27><12>  ( .D(n18487), .E(n18421), .CK(clk), .Q(
        \RAM<27><12> ) );
  EDFFX1 \RAM_reg<27><11>  ( .D(n18483), .E(n18421), .CK(clk), .Q(
        \RAM<27><11> ) );
  EDFFX1 \RAM_reg<27><10>  ( .D(n18479), .E(n18421), .CK(clk), .Q(
        \RAM<27><10> ) );
  EDFFX1 \RAM_reg<27><9>  ( .D(n18475), .E(n18421), .CK(clk), .Q(\RAM<27><9> )
         );
  EDFFX1 \RAM_reg<27><8>  ( .D(n18471), .E(n18421), .CK(clk), .Q(\RAM<27><8> )
         );
  EDFFX1 \RAM_reg<27><7>  ( .D(n18467), .E(n3523), .CK(clk), .Q(\RAM<27><7> )
         );
  EDFFX1 \RAM_reg<27><6>  ( .D(n18463), .E(n3523), .CK(clk), .Q(\RAM<27><6> )
         );
  EDFFX1 \RAM_reg<27><5>  ( .D(n18459), .E(n18420), .CK(clk), .Q(\RAM<27><5> )
         );
  EDFFX1 \RAM_reg<27><4>  ( .D(n18455), .E(n18421), .CK(clk), .Q(\RAM<27><4> )
         );
  EDFFX1 \RAM_reg<27><3>  ( .D(n18451), .E(n18420), .CK(clk), .Q(\RAM<27><3> )
         );
  EDFFX1 \RAM_reg<27><2>  ( .D(n18447), .E(n18421), .CK(clk), .Q(\RAM<27><2> )
         );
  EDFFX1 \RAM_reg<27><1>  ( .D(n18443), .E(n18420), .CK(clk), .Q(\RAM<27><1> )
         );
  EDFFX1 \RAM_reg<27><0>  ( .D(n18439), .E(n18421), .CK(clk), .Q(\RAM<27><0> )
         );
  EDFFX1 \RAM_reg<23><31>  ( .D(n18563), .E(n18312), .CK(clk), .Q(
        \RAM<23><31> ) );
  EDFFX1 \RAM_reg<23><30>  ( .D(n18559), .E(n18312), .CK(clk), .Q(
        \RAM<23><30> ) );
  EDFFX1 \RAM_reg<23><29>  ( .D(n18555), .E(n18312), .CK(clk), .Q(
        \RAM<23><29> ) );
  EDFFX1 \RAM_reg<23><28>  ( .D(n18551), .E(n18312), .CK(clk), .Q(
        \RAM<23><28> ) );
  EDFFX1 \RAM_reg<23><27>  ( .D(n18547), .E(n18312), .CK(clk), .Q(
        \RAM<23><27> ) );
  EDFFX1 \RAM_reg<23><26>  ( .D(n18543), .E(n18312), .CK(clk), .Q(
        \RAM<23><26> ) );
  EDFFX1 \RAM_reg<23><25>  ( .D(n18539), .E(n18312), .CK(clk), .Q(
        \RAM<23><25> ) );
  EDFFX1 \RAM_reg<23><24>  ( .D(n18535), .E(n18312), .CK(clk), .Q(
        \RAM<23><24> ) );
  EDFFX1 \RAM_reg<23><23>  ( .D(n18531), .E(n18312), .CK(clk), .Q(
        \RAM<23><23> ) );
  EDFFX1 \RAM_reg<23><22>  ( .D(n18527), .E(n18312), .CK(clk), .Q(
        \RAM<23><22> ) );
  EDFFX1 \RAM_reg<23><21>  ( .D(n18523), .E(n18312), .CK(clk), .Q(
        \RAM<23><21> ) );
  EDFFX1 \RAM_reg<23><20>  ( .D(n18519), .E(n18312), .CK(clk), .Q(
        \RAM<23><20> ) );
  EDFFX1 \RAM_reg<23><19>  ( .D(n18515), .E(n18313), .CK(clk), .Q(
        \RAM<23><19> ) );
  EDFFX1 \RAM_reg<23><18>  ( .D(n18511), .E(n18313), .CK(clk), .Q(
        \RAM<23><18> ) );
  EDFFX1 \RAM_reg<23><17>  ( .D(n18507), .E(n18313), .CK(clk), .Q(
        \RAM<23><17> ) );
  EDFFX1 \RAM_reg<23><16>  ( .D(n18503), .E(n18313), .CK(clk), .Q(
        \RAM<23><16> ) );
  EDFFX1 \RAM_reg<23><15>  ( .D(n18499), .E(n18313), .CK(clk), .Q(
        \RAM<23><15> ) );
  EDFFX1 \RAM_reg<23><14>  ( .D(n18495), .E(n18313), .CK(clk), .Q(
        \RAM<23><14> ) );
  EDFFX1 \RAM_reg<23><13>  ( .D(n18491), .E(n18313), .CK(clk), .Q(
        \RAM<23><13> ) );
  EDFFX1 \RAM_reg<23><12>  ( .D(n18487), .E(n18313), .CK(clk), .Q(
        \RAM<23><12> ) );
  EDFFX1 \RAM_reg<23><11>  ( .D(n18483), .E(n18313), .CK(clk), .Q(
        \RAM<23><11> ) );
  EDFFX1 \RAM_reg<23><10>  ( .D(n18479), .E(n18313), .CK(clk), .Q(
        \RAM<23><10> ) );
  EDFFX1 \RAM_reg<23><9>  ( .D(n18475), .E(n18313), .CK(clk), .Q(\RAM<23><9> )
         );
  EDFFX1 \RAM_reg<23><8>  ( .D(n18471), .E(n18313), .CK(clk), .Q(\RAM<23><8> )
         );
  EDFFX1 \RAM_reg<23><7>  ( .D(n18467), .E(n3563), .CK(clk), .Q(\RAM<23><7> )
         );
  EDFFX1 \RAM_reg<23><6>  ( .D(n18463), .E(n3563), .CK(clk), .Q(\RAM<23><6> )
         );
  EDFFX1 \RAM_reg<23><5>  ( .D(n18459), .E(n18312), .CK(clk), .Q(\RAM<23><5> )
         );
  EDFFX1 \RAM_reg<23><4>  ( .D(n18455), .E(n18313), .CK(clk), .Q(\RAM<23><4> )
         );
  EDFFX1 \RAM_reg<23><3>  ( .D(n18451), .E(n18312), .CK(clk), .Q(\RAM<23><3> )
         );
  EDFFX1 \RAM_reg<23><2>  ( .D(n18447), .E(n18313), .CK(clk), .Q(\RAM<23><2> )
         );
  EDFFX1 \RAM_reg<23><1>  ( .D(n18443), .E(n18312), .CK(clk), .Q(\RAM<23><1> )
         );
  EDFFX1 \RAM_reg<23><0>  ( .D(n18439), .E(n18313), .CK(clk), .Q(\RAM<23><0> )
         );
  EDFFX1 \RAM_reg<19><31>  ( .D(n18563), .E(n18423), .CK(clk), .Q(
        \RAM<19><31> ) );
  EDFFX1 \RAM_reg<19><30>  ( .D(n18559), .E(n18423), .CK(clk), .Q(
        \RAM<19><30> ) );
  EDFFX1 \RAM_reg<19><29>  ( .D(n18555), .E(n18423), .CK(clk), .Q(
        \RAM<19><29> ) );
  EDFFX1 \RAM_reg<19><28>  ( .D(n18551), .E(n18423), .CK(clk), .Q(
        \RAM<19><28> ) );
  EDFFX1 \RAM_reg<19><27>  ( .D(n18547), .E(n18423), .CK(clk), .Q(
        \RAM<19><27> ) );
  EDFFX1 \RAM_reg<19><26>  ( .D(n18543), .E(n18423), .CK(clk), .Q(
        \RAM<19><26> ) );
  EDFFX1 \RAM_reg<19><25>  ( .D(n18539), .E(n18423), .CK(clk), .Q(
        \RAM<19><25> ) );
  EDFFX1 \RAM_reg<19><24>  ( .D(n18535), .E(n18423), .CK(clk), .Q(
        \RAM<19><24> ) );
  EDFFX1 \RAM_reg<19><23>  ( .D(n18531), .E(n18423), .CK(clk), .Q(
        \RAM<19><23> ) );
  EDFFX1 \RAM_reg<19><22>  ( .D(n18527), .E(n18423), .CK(clk), .Q(
        \RAM<19><22> ) );
  EDFFX1 \RAM_reg<19><21>  ( .D(n18523), .E(n18423), .CK(clk), .Q(
        \RAM<19><21> ) );
  EDFFX1 \RAM_reg<19><20>  ( .D(n18519), .E(n18423), .CK(clk), .Q(
        \RAM<19><20> ) );
  EDFFX1 \RAM_reg<19><19>  ( .D(n18515), .E(n18424), .CK(clk), .Q(
        \RAM<19><19> ) );
  EDFFX1 \RAM_reg<19><18>  ( .D(n18511), .E(n18424), .CK(clk), .Q(
        \RAM<19><18> ) );
  EDFFX1 \RAM_reg<19><17>  ( .D(n18507), .E(n18424), .CK(clk), .Q(
        \RAM<19><17> ) );
  EDFFX1 \RAM_reg<19><16>  ( .D(n18503), .E(n18424), .CK(clk), .Q(
        \RAM<19><16> ) );
  EDFFX1 \RAM_reg<19><15>  ( .D(n18499), .E(n18424), .CK(clk), .Q(
        \RAM<19><15> ) );
  EDFFX1 \RAM_reg<19><14>  ( .D(n18495), .E(n18424), .CK(clk), .Q(
        \RAM<19><14> ) );
  EDFFX1 \RAM_reg<19><13>  ( .D(n18491), .E(n18424), .CK(clk), .Q(
        \RAM<19><13> ) );
  EDFFX1 \RAM_reg<19><12>  ( .D(n18487), .E(n18424), .CK(clk), .Q(
        \RAM<19><12> ) );
  EDFFX1 \RAM_reg<19><11>  ( .D(n18483), .E(n18424), .CK(clk), .Q(
        \RAM<19><11> ) );
  EDFFX1 \RAM_reg<19><10>  ( .D(n18479), .E(n18424), .CK(clk), .Q(
        \RAM<19><10> ) );
  EDFFX1 \RAM_reg<19><9>  ( .D(n18475), .E(n18424), .CK(clk), .Q(\RAM<19><9> )
         );
  EDFFX1 \RAM_reg<19><8>  ( .D(n18471), .E(n18424), .CK(clk), .Q(\RAM<19><8> )
         );
  EDFFX1 \RAM_reg<19><7>  ( .D(n18467), .E(n3522), .CK(clk), .Q(\RAM<19><7> )
         );
  EDFFX1 \RAM_reg<19><6>  ( .D(n18463), .E(n3522), .CK(clk), .Q(\RAM<19><6> )
         );
  EDFFX1 \RAM_reg<19><5>  ( .D(n18459), .E(n18423), .CK(clk), .Q(\RAM<19><5> )
         );
  EDFFX1 \RAM_reg<19><4>  ( .D(n18455), .E(n18424), .CK(clk), .Q(\RAM<19><4> )
         );
  EDFFX1 \RAM_reg<19><3>  ( .D(n18451), .E(n18423), .CK(clk), .Q(\RAM<19><3> )
         );
  EDFFX1 \RAM_reg<19><2>  ( .D(n18447), .E(n18424), .CK(clk), .Q(\RAM<19><2> )
         );
  EDFFX1 \RAM_reg<19><1>  ( .D(n18443), .E(n18423), .CK(clk), .Q(\RAM<19><1> )
         );
  EDFFX1 \RAM_reg<19><0>  ( .D(n18439), .E(n18424), .CK(clk), .Q(\RAM<19><0> )
         );
  EDFFX1 \RAM_reg<15><31>  ( .D(n18563), .E(n18318), .CK(clk), .Q(
        \RAM<15><31> ) );
  EDFFX1 \RAM_reg<15><30>  ( .D(n18559), .E(n18318), .CK(clk), .Q(
        \RAM<15><30> ) );
  EDFFX1 \RAM_reg<15><29>  ( .D(n18555), .E(n18318), .CK(clk), .Q(
        \RAM<15><29> ) );
  EDFFX1 \RAM_reg<15><28>  ( .D(n18551), .E(n18318), .CK(clk), .Q(
        \RAM<15><28> ) );
  EDFFX1 \RAM_reg<15><27>  ( .D(n18547), .E(n18318), .CK(clk), .Q(
        \RAM<15><27> ) );
  EDFFX1 \RAM_reg<15><26>  ( .D(n18543), .E(n18318), .CK(clk), .Q(
        \RAM<15><26> ) );
  EDFFX1 \RAM_reg<15><25>  ( .D(n18539), .E(n18318), .CK(clk), .Q(
        \RAM<15><25> ) );
  EDFFX1 \RAM_reg<15><24>  ( .D(n18535), .E(n18318), .CK(clk), .Q(
        \RAM<15><24> ) );
  EDFFX1 \RAM_reg<15><23>  ( .D(n18531), .E(n18318), .CK(clk), .Q(
        \RAM<15><23> ) );
  EDFFX1 \RAM_reg<15><22>  ( .D(n18527), .E(n18318), .CK(clk), .Q(
        \RAM<15><22> ) );
  EDFFX1 \RAM_reg<15><21>  ( .D(n18523), .E(n18318), .CK(clk), .Q(
        \RAM<15><21> ) );
  EDFFX1 \RAM_reg<15><20>  ( .D(n18519), .E(n18318), .CK(clk), .Q(
        \RAM<15><20> ) );
  EDFFX1 \RAM_reg<15><19>  ( .D(n18515), .E(n18319), .CK(clk), .Q(
        \RAM<15><19> ) );
  EDFFX1 \RAM_reg<15><18>  ( .D(n18511), .E(n18319), .CK(clk), .Q(
        \RAM<15><18> ) );
  EDFFX1 \RAM_reg<15><17>  ( .D(n18507), .E(n18319), .CK(clk), .Q(
        \RAM<15><17> ) );
  EDFFX1 \RAM_reg<15><16>  ( .D(n18503), .E(n18319), .CK(clk), .Q(
        \RAM<15><16> ) );
  EDFFX1 \RAM_reg<15><15>  ( .D(n18499), .E(n18319), .CK(clk), .Q(
        \RAM<15><15> ) );
  EDFFX1 \RAM_reg<15><14>  ( .D(n18495), .E(n18319), .CK(clk), .Q(
        \RAM<15><14> ) );
  EDFFX1 \RAM_reg<15><13>  ( .D(n18491), .E(n18319), .CK(clk), .Q(
        \RAM<15><13> ) );
  EDFFX1 \RAM_reg<15><12>  ( .D(n18487), .E(n18319), .CK(clk), .Q(
        \RAM<15><12> ) );
  EDFFX1 \RAM_reg<15><11>  ( .D(n18483), .E(n18319), .CK(clk), .Q(
        \RAM<15><11> ) );
  EDFFX1 \RAM_reg<15><10>  ( .D(n18479), .E(n18319), .CK(clk), .Q(
        \RAM<15><10> ) );
  EDFFX1 \RAM_reg<15><9>  ( .D(n18475), .E(n18319), .CK(clk), .Q(\RAM<15><9> )
         );
  EDFFX1 \RAM_reg<15><8>  ( .D(n18471), .E(n18319), .CK(clk), .Q(\RAM<15><8> )
         );
  EDFFX1 \RAM_reg<15><7>  ( .D(n18467), .E(n3559), .CK(clk), .Q(\RAM<15><7> )
         );
  EDFFX1 \RAM_reg<15><6>  ( .D(n18463), .E(n3559), .CK(clk), .Q(\RAM<15><6> )
         );
  EDFFX1 \RAM_reg<15><5>  ( .D(n18459), .E(n18318), .CK(clk), .Q(\RAM<15><5> )
         );
  EDFFX1 \RAM_reg<15><4>  ( .D(n18455), .E(n18319), .CK(clk), .Q(\RAM<15><4> )
         );
  EDFFX1 \RAM_reg<15><3>  ( .D(n18451), .E(n18318), .CK(clk), .Q(\RAM<15><3> )
         );
  EDFFX1 \RAM_reg<15><2>  ( .D(n18447), .E(n18319), .CK(clk), .Q(\RAM<15><2> )
         );
  EDFFX1 \RAM_reg<15><1>  ( .D(n18443), .E(n18318), .CK(clk), .Q(\RAM<15><1> )
         );
  EDFFX1 \RAM_reg<15><0>  ( .D(n18439), .E(n18319), .CK(clk), .Q(\RAM<15><0> )
         );
  EDFFX1 \RAM_reg<11><31>  ( .D(n18563), .E(n18282), .CK(clk), .Q(
        \RAM<11><31> ) );
  EDFFX1 \RAM_reg<11><30>  ( .D(n18559), .E(n18282), .CK(clk), .Q(
        \RAM<11><30> ) );
  EDFFX1 \RAM_reg<11><29>  ( .D(n18555), .E(n18282), .CK(clk), .Q(
        \RAM<11><29> ) );
  EDFFX1 \RAM_reg<11><28>  ( .D(n18551), .E(n18282), .CK(clk), .Q(
        \RAM<11><28> ) );
  EDFFX1 \RAM_reg<11><27>  ( .D(n18547), .E(n18282), .CK(clk), .Q(
        \RAM<11><27> ) );
  EDFFX1 \RAM_reg<11><26>  ( .D(n18543), .E(n18282), .CK(clk), .Q(
        \RAM<11><26> ) );
  EDFFX1 \RAM_reg<11><25>  ( .D(n18539), .E(n18282), .CK(clk), .Q(
        \RAM<11><25> ) );
  EDFFX1 \RAM_reg<11><24>  ( .D(n18535), .E(n18282), .CK(clk), .Q(
        \RAM<11><24> ) );
  EDFFX1 \RAM_reg<11><23>  ( .D(n18531), .E(n18282), .CK(clk), .Q(
        \RAM<11><23> ) );
  EDFFX1 \RAM_reg<11><22>  ( .D(n18527), .E(n18282), .CK(clk), .Q(
        \RAM<11><22> ) );
  EDFFX1 \RAM_reg<11><21>  ( .D(n18523), .E(n18282), .CK(clk), .Q(
        \RAM<11><21> ) );
  EDFFX1 \RAM_reg<11><20>  ( .D(n18519), .E(n18282), .CK(clk), .Q(
        \RAM<11><20> ) );
  EDFFX1 \RAM_reg<11><19>  ( .D(n18515), .E(n18283), .CK(clk), .Q(
        \RAM<11><19> ) );
  EDFFX1 \RAM_reg<11><18>  ( .D(n18511), .E(n18283), .CK(clk), .Q(
        \RAM<11><18> ) );
  EDFFX1 \RAM_reg<11><17>  ( .D(n18507), .E(n18283), .CK(clk), .Q(
        \RAM<11><17> ) );
  EDFFX1 \RAM_reg<11><16>  ( .D(n18503), .E(n18283), .CK(clk), .Q(
        \RAM<11><16> ) );
  EDFFX1 \RAM_reg<11><15>  ( .D(n18499), .E(n18283), .CK(clk), .Q(
        \RAM<11><15> ) );
  EDFFX1 \RAM_reg<11><14>  ( .D(n18495), .E(n18283), .CK(clk), .Q(
        \RAM<11><14> ) );
  EDFFX1 \RAM_reg<11><13>  ( .D(n18491), .E(n18283), .CK(clk), .Q(
        \RAM<11><13> ) );
  EDFFX1 \RAM_reg<11><12>  ( .D(n18487), .E(n18283), .CK(clk), .Q(
        \RAM<11><12> ) );
  EDFFX1 \RAM_reg<11><11>  ( .D(n18483), .E(n18283), .CK(clk), .Q(
        \RAM<11><11> ) );
  EDFFX1 \RAM_reg<11><10>  ( .D(n18479), .E(n18283), .CK(clk), .Q(
        \RAM<11><10> ) );
  EDFFX1 \RAM_reg<11><9>  ( .D(n18475), .E(n18283), .CK(clk), .Q(\RAM<11><9> )
         );
  EDFFX1 \RAM_reg<11><8>  ( .D(n18471), .E(n18283), .CK(clk), .Q(\RAM<11><8> )
         );
  EDFFX1 \RAM_reg<11><7>  ( .D(n18467), .E(n3577), .CK(clk), .Q(\RAM<11><7> )
         );
  EDFFX1 \RAM_reg<11><6>  ( .D(n18463), .E(n3577), .CK(clk), .Q(\RAM<11><6> )
         );
  EDFFX1 \RAM_reg<11><5>  ( .D(n18459), .E(n18282), .CK(clk), .Q(\RAM<11><5> )
         );
  EDFFX1 \RAM_reg<11><4>  ( .D(n18455), .E(n18283), .CK(clk), .Q(\RAM<11><4> )
         );
  EDFFX1 \RAM_reg<11><3>  ( .D(n18451), .E(n18282), .CK(clk), .Q(\RAM<11><3> )
         );
  EDFFX1 \RAM_reg<11><2>  ( .D(n18447), .E(n18283), .CK(clk), .Q(\RAM<11><2> )
         );
  EDFFX1 \RAM_reg<11><1>  ( .D(n18443), .E(n18282), .CK(clk), .Q(\RAM<11><1> )
         );
  EDFFX1 \RAM_reg<11><0>  ( .D(n18439), .E(n18283), .CK(clk), .Q(\RAM<11><0> )
         );
  EDFFX1 \RAM_reg<7><31>  ( .D(n18563), .E(n18435), .CK(clk), .Q(\RAM<7><31> )
         );
  EDFFX1 \RAM_reg<7><30>  ( .D(n18559), .E(n18435), .CK(clk), .Q(\RAM<7><30> )
         );
  EDFFX1 \RAM_reg<7><29>  ( .D(n18555), .E(n18435), .CK(clk), .Q(\RAM<7><29> )
         );
  EDFFX1 \RAM_reg<7><28>  ( .D(n18551), .E(n18435), .CK(clk), .Q(\RAM<7><28> )
         );
  EDFFX1 \RAM_reg<7><27>  ( .D(n18547), .E(n18435), .CK(clk), .Q(\RAM<7><27> )
         );
  EDFFX1 \RAM_reg<7><26>  ( .D(n18543), .E(n18435), .CK(clk), .Q(\RAM<7><26> )
         );
  EDFFX1 \RAM_reg<7><25>  ( .D(n18539), .E(n18435), .CK(clk), .Q(\RAM<7><25> )
         );
  EDFFX1 \RAM_reg<7><24>  ( .D(n18535), .E(n18435), .CK(clk), .Q(\RAM<7><24> )
         );
  EDFFX1 \RAM_reg<7><23>  ( .D(n18531), .E(n18435), .CK(clk), .Q(\RAM<7><23> )
         );
  EDFFX1 \RAM_reg<7><22>  ( .D(n18527), .E(n18435), .CK(clk), .Q(\RAM<7><22> )
         );
  EDFFX1 \RAM_reg<7><21>  ( .D(n18523), .E(n18435), .CK(clk), .Q(\RAM<7><21> )
         );
  EDFFX1 \RAM_reg<7><20>  ( .D(n18519), .E(n18435), .CK(clk), .Q(\RAM<7><20> )
         );
  EDFFX1 \RAM_reg<7><19>  ( .D(n18515), .E(n18436), .CK(clk), .Q(\RAM<7><19> )
         );
  EDFFX1 \RAM_reg<7><18>  ( .D(n18511), .E(n18436), .CK(clk), .Q(\RAM<7><18> )
         );
  EDFFX1 \RAM_reg<7><17>  ( .D(n18507), .E(n18436), .CK(clk), .Q(\RAM<7><17> )
         );
  EDFFX1 \RAM_reg<7><16>  ( .D(n18503), .E(n18436), .CK(clk), .Q(\RAM<7><16> )
         );
  EDFFX1 \RAM_reg<7><15>  ( .D(n18499), .E(n18436), .CK(clk), .Q(\RAM<7><15> )
         );
  EDFFX1 \RAM_reg<7><14>  ( .D(n18495), .E(n18436), .CK(clk), .Q(\RAM<7><14> )
         );
  EDFFX1 \RAM_reg<7><13>  ( .D(n18491), .E(n18436), .CK(clk), .Q(\RAM<7><13> )
         );
  EDFFX1 \RAM_reg<7><12>  ( .D(n18487), .E(n18436), .CK(clk), .Q(\RAM<7><12> )
         );
  EDFFX1 \RAM_reg<7><11>  ( .D(n18483), .E(n18436), .CK(clk), .Q(\RAM<7><11> )
         );
  EDFFX1 \RAM_reg<7><10>  ( .D(n18479), .E(n18436), .CK(clk), .Q(\RAM<7><10> )
         );
  EDFFX1 \RAM_reg<7><9>  ( .D(n18475), .E(n18436), .CK(clk), .Q(\RAM<7><9> )
         );
  EDFFX1 \RAM_reg<7><8>  ( .D(n18471), .E(n18436), .CK(clk), .Q(\RAM<7><8> )
         );
  EDFFX1 \RAM_reg<7><7>  ( .D(n18467), .E(n66), .CK(clk), .Q(\RAM<7><7> ) );
  EDFFX1 \RAM_reg<7><6>  ( .D(n18463), .E(n66), .CK(clk), .Q(\RAM<7><6> ) );
  EDFFX1 \RAM_reg<7><5>  ( .D(n18459), .E(n18435), .CK(clk), .Q(\RAM<7><5> )
         );
  EDFFX1 \RAM_reg<7><4>  ( .D(n18455), .E(n18436), .CK(clk), .Q(\RAM<7><4> )
         );
  EDFFX1 \RAM_reg<7><3>  ( .D(n18451), .E(n18435), .CK(clk), .Q(\RAM<7><3> )
         );
  EDFFX1 \RAM_reg<7><2>  ( .D(n18447), .E(n18436), .CK(clk), .Q(\RAM<7><2> )
         );
  EDFFX1 \RAM_reg<7><1>  ( .D(n18443), .E(n18435), .CK(clk), .Q(\RAM<7><1> )
         );
  EDFFX1 \RAM_reg<7><0>  ( .D(n18439), .E(n18436), .CK(clk), .Q(\RAM<7><0> )
         );
  EDFFX1 \RAM_reg<3><31>  ( .D(n18563), .E(n18288), .CK(clk), .Q(\RAM<3><31> )
         );
  EDFFX1 \RAM_reg<3><30>  ( .D(n18559), .E(n18288), .CK(clk), .Q(\RAM<3><30> )
         );
  EDFFX1 \RAM_reg<3><29>  ( .D(n18555), .E(n18288), .CK(clk), .Q(\RAM<3><29> )
         );
  EDFFX1 \RAM_reg<3><28>  ( .D(n18551), .E(n18288), .CK(clk), .Q(\RAM<3><28> )
         );
  EDFFX1 \RAM_reg<3><27>  ( .D(n18547), .E(n18288), .CK(clk), .Q(\RAM<3><27> )
         );
  EDFFX1 \RAM_reg<3><26>  ( .D(n18543), .E(n18288), .CK(clk), .Q(\RAM<3><26> )
         );
  EDFFX1 \RAM_reg<3><25>  ( .D(n18539), .E(n18288), .CK(clk), .Q(\RAM<3><25> )
         );
  EDFFX1 \RAM_reg<3><24>  ( .D(n18535), .E(n18288), .CK(clk), .Q(\RAM<3><24> )
         );
  EDFFX1 \RAM_reg<3><23>  ( .D(n18531), .E(n18288), .CK(clk), .Q(\RAM<3><23> )
         );
  EDFFX1 \RAM_reg<3><22>  ( .D(n18527), .E(n18288), .CK(clk), .Q(\RAM<3><22> )
         );
  EDFFX1 \RAM_reg<3><21>  ( .D(n18523), .E(n18288), .CK(clk), .Q(\RAM<3><21> )
         );
  EDFFX1 \RAM_reg<3><20>  ( .D(n18519), .E(n18288), .CK(clk), .Q(\RAM<3><20> )
         );
  EDFFX1 \RAM_reg<3><19>  ( .D(n18515), .E(n18289), .CK(clk), .Q(\RAM<3><19> )
         );
  EDFFX1 \RAM_reg<3><18>  ( .D(n18511), .E(n18289), .CK(clk), .Q(\RAM<3><18> )
         );
  EDFFX1 \RAM_reg<3><17>  ( .D(n18507), .E(n18289), .CK(clk), .Q(\RAM<3><17> )
         );
  EDFFX1 \RAM_reg<3><16>  ( .D(n18503), .E(n18289), .CK(clk), .Q(\RAM<3><16> )
         );
  EDFFX1 \RAM_reg<3><15>  ( .D(n18499), .E(n18289), .CK(clk), .Q(\RAM<3><15> )
         );
  EDFFX1 \RAM_reg<3><14>  ( .D(n18495), .E(n18289), .CK(clk), .Q(\RAM<3><14> )
         );
  EDFFX1 \RAM_reg<3><13>  ( .D(n18491), .E(n18289), .CK(clk), .Q(\RAM<3><13> )
         );
  EDFFX1 \RAM_reg<3><12>  ( .D(n18487), .E(n18289), .CK(clk), .Q(\RAM<3><12> )
         );
  EDFFX1 \RAM_reg<3><11>  ( .D(n18483), .E(n18289), .CK(clk), .Q(\RAM<3><11> )
         );
  EDFFX1 \RAM_reg<3><10>  ( .D(n18479), .E(n18289), .CK(clk), .Q(\RAM<3><10> )
         );
  EDFFX1 \RAM_reg<3><9>  ( .D(n18475), .E(n18289), .CK(clk), .Q(\RAM<3><9> )
         );
  EDFFX1 \RAM_reg<3><8>  ( .D(n18471), .E(n18289), .CK(clk), .Q(\RAM<3><8> )
         );
  EDFFX1 \RAM_reg<3><7>  ( .D(n18467), .E(n3574), .CK(clk), .Q(\RAM<3><7> ) );
  EDFFX1 \RAM_reg<3><6>  ( .D(n18463), .E(n3574), .CK(clk), .Q(\RAM<3><6> ) );
  EDFFX1 \RAM_reg<3><5>  ( .D(n18459), .E(n18288), .CK(clk), .Q(\RAM<3><5> )
         );
  EDFFX1 \RAM_reg<3><4>  ( .D(n18455), .E(n18289), .CK(clk), .Q(\RAM<3><4> )
         );
  EDFFX1 \RAM_reg<3><3>  ( .D(n18451), .E(n18288), .CK(clk), .Q(\RAM<3><3> )
         );
  EDFFX1 \RAM_reg<3><2>  ( .D(n18447), .E(n18289), .CK(clk), .Q(\RAM<3><2> )
         );
  EDFFX1 \RAM_reg<3><1>  ( .D(n18443), .E(n18288), .CK(clk), .Q(\RAM<3><1> )
         );
  EDFFX1 \RAM_reg<3><0>  ( .D(n18439), .E(n18289), .CK(clk), .Q(\RAM<3><0> )
         );
  EDFFX1 \RAM_reg<58><31>  ( .D(\wd<31> ), .E(n18330), .CK(clk), .Q(
        \RAM<58><31> ) );
  EDFFX1 \RAM_reg<58><30>  ( .D(\wd<30> ), .E(n18330), .CK(clk), .Q(
        \RAM<58><30> ) );
  EDFFX1 \RAM_reg<58><29>  ( .D(\wd<29> ), .E(n18330), .CK(clk), .Q(
        \RAM<58><29> ) );
  EDFFX1 \RAM_reg<58><28>  ( .D(\wd<28> ), .E(n18330), .CK(clk), .Q(
        \RAM<58><28> ) );
  EDFFX1 \RAM_reg<58><27>  ( .D(\wd<27> ), .E(n18330), .CK(clk), .Q(
        \RAM<58><27> ) );
  EDFFX1 \RAM_reg<58><26>  ( .D(\wd<26> ), .E(n18330), .CK(clk), .Q(
        \RAM<58><26> ) );
  EDFFX1 \RAM_reg<58><25>  ( .D(\wd<25> ), .E(n18330), .CK(clk), .Q(
        \RAM<58><25> ) );
  EDFFX1 \RAM_reg<58><24>  ( .D(\wd<24> ), .E(n18330), .CK(clk), .Q(
        \RAM<58><24> ) );
  EDFFX1 \RAM_reg<58><23>  ( .D(\wd<23> ), .E(n18330), .CK(clk), .Q(
        \RAM<58><23> ) );
  EDFFX1 \RAM_reg<58><22>  ( .D(\wd<22> ), .E(n18330), .CK(clk), .Q(
        \RAM<58><22> ) );
  EDFFX1 \RAM_reg<58><21>  ( .D(\wd<21> ), .E(n18330), .CK(clk), .Q(
        \RAM<58><21> ) );
  EDFFX1 \RAM_reg<58><20>  ( .D(\wd<20> ), .E(n18330), .CK(clk), .Q(
        \RAM<58><20> ) );
  EDFFX1 \RAM_reg<58><19>  ( .D(\wd<19> ), .E(n18331), .CK(clk), .Q(
        \RAM<58><19> ) );
  EDFFX1 \RAM_reg<58><18>  ( .D(\wd<18> ), .E(n18331), .CK(clk), .Q(
        \RAM<58><18> ) );
  EDFFX1 \RAM_reg<58><17>  ( .D(\wd<17> ), .E(n18331), .CK(clk), .Q(
        \RAM<58><17> ) );
  EDFFX1 \RAM_reg<58><16>  ( .D(\wd<16> ), .E(n18331), .CK(clk), .Q(
        \RAM<58><16> ) );
  EDFFX1 \RAM_reg<58><15>  ( .D(\wd<15> ), .E(n18331), .CK(clk), .Q(
        \RAM<58><15> ) );
  EDFFX1 \RAM_reg<58><14>  ( .D(\wd<14> ), .E(n18331), .CK(clk), .Q(
        \RAM<58><14> ) );
  EDFFX1 \RAM_reg<58><13>  ( .D(\wd<13> ), .E(n18331), .CK(clk), .Q(
        \RAM<58><13> ) );
  EDFFX1 \RAM_reg<58><12>  ( .D(\wd<12> ), .E(n18331), .CK(clk), .Q(
        \RAM<58><12> ) );
  EDFFX1 \RAM_reg<58><11>  ( .D(\wd<11> ), .E(n18331), .CK(clk), .Q(
        \RAM<58><11> ) );
  EDFFX1 \RAM_reg<58><10>  ( .D(\wd<10> ), .E(n18331), .CK(clk), .Q(
        \RAM<58><10> ) );
  EDFFX1 \RAM_reg<58><9>  ( .D(\wd<9> ), .E(n18331), .CK(clk), .Q(\RAM<58><9> ) );
  EDFFX1 \RAM_reg<58><8>  ( .D(\wd<8> ), .E(n18331), .CK(clk), .Q(\RAM<58><8> ) );
  EDFFX1 \RAM_reg<58><7>  ( .D(\wd<7> ), .E(n3555), .CK(clk), .Q(\RAM<58><7> )
         );
  EDFFX1 \RAM_reg<58><6>  ( .D(\wd<6> ), .E(n3555), .CK(clk), .Q(\RAM<58><6> )
         );
  EDFFX1 \RAM_reg<58><5>  ( .D(\wd<5> ), .E(n18330), .CK(clk), .Q(\RAM<58><5> ) );
  EDFFX1 \RAM_reg<58><4>  ( .D(\wd<4> ), .E(n18331), .CK(clk), .Q(\RAM<58><4> ) );
  EDFFX1 \RAM_reg<58><3>  ( .D(\wd<3> ), .E(n18330), .CK(clk), .Q(\RAM<58><3> ) );
  EDFFX1 \RAM_reg<58><2>  ( .D(\wd<2> ), .E(n18331), .CK(clk), .Q(\RAM<58><2> ) );
  EDFFX1 \RAM_reg<58><1>  ( .D(\wd<1> ), .E(n18330), .CK(clk), .Q(\RAM<58><1> ) );
  EDFFX1 \RAM_reg<58><0>  ( .D(\wd<0> ), .E(n18331), .CK(clk), .Q(\RAM<58><0> ) );
  EDFFX1 \RAM_reg<50><31>  ( .D(\wd<31> ), .E(n18336), .CK(clk), .Q(
        \RAM<50><31> ) );
  EDFFX1 \RAM_reg<50><30>  ( .D(\wd<30> ), .E(n18336), .CK(clk), .Q(
        \RAM<50><30> ) );
  EDFFX1 \RAM_reg<50><29>  ( .D(\wd<29> ), .E(n18336), .CK(clk), .Q(
        \RAM<50><29> ) );
  EDFFX1 \RAM_reg<50><28>  ( .D(\wd<28> ), .E(n18336), .CK(clk), .Q(
        \RAM<50><28> ) );
  EDFFX1 \RAM_reg<50><27>  ( .D(\wd<27> ), .E(n18336), .CK(clk), .Q(
        \RAM<50><27> ) );
  EDFFX1 \RAM_reg<50><26>  ( .D(\wd<26> ), .E(n18336), .CK(clk), .Q(
        \RAM<50><26> ) );
  EDFFX1 \RAM_reg<50><25>  ( .D(\wd<25> ), .E(n18336), .CK(clk), .Q(
        \RAM<50><25> ) );
  EDFFX1 \RAM_reg<50><24>  ( .D(\wd<24> ), .E(n18336), .CK(clk), .Q(
        \RAM<50><24> ) );
  EDFFX1 \RAM_reg<50><23>  ( .D(\wd<23> ), .E(n18336), .CK(clk), .Q(
        \RAM<50><23> ) );
  EDFFX1 \RAM_reg<50><22>  ( .D(\wd<22> ), .E(n18336), .CK(clk), .Q(
        \RAM<50><22> ) );
  EDFFX1 \RAM_reg<50><21>  ( .D(\wd<21> ), .E(n18336), .CK(clk), .Q(
        \RAM<50><21> ) );
  EDFFX1 \RAM_reg<50><20>  ( .D(\wd<20> ), .E(n18336), .CK(clk), .Q(
        \RAM<50><20> ) );
  EDFFX1 \RAM_reg<50><19>  ( .D(\wd<19> ), .E(n18337), .CK(clk), .Q(
        \RAM<50><19> ) );
  EDFFX1 \RAM_reg<50><18>  ( .D(\wd<18> ), .E(n18337), .CK(clk), .Q(
        \RAM<50><18> ) );
  EDFFX1 \RAM_reg<50><17>  ( .D(\wd<17> ), .E(n18337), .CK(clk), .Q(
        \RAM<50><17> ) );
  EDFFX1 \RAM_reg<50><16>  ( .D(\wd<16> ), .E(n18337), .CK(clk), .Q(
        \RAM<50><16> ) );
  EDFFX1 \RAM_reg<50><15>  ( .D(\wd<15> ), .E(n18337), .CK(clk), .Q(
        \RAM<50><15> ) );
  EDFFX1 \RAM_reg<50><14>  ( .D(\wd<14> ), .E(n18337), .CK(clk), .Q(
        \RAM<50><14> ) );
  EDFFX1 \RAM_reg<50><13>  ( .D(\wd<13> ), .E(n18337), .CK(clk), .Q(
        \RAM<50><13> ) );
  EDFFX1 \RAM_reg<50><12>  ( .D(\wd<12> ), .E(n18337), .CK(clk), .Q(
        \RAM<50><12> ) );
  EDFFX1 \RAM_reg<50><11>  ( .D(\wd<11> ), .E(n18337), .CK(clk), .Q(
        \RAM<50><11> ) );
  EDFFX1 \RAM_reg<50><10>  ( .D(\wd<10> ), .E(n18337), .CK(clk), .Q(
        \RAM<50><10> ) );
  EDFFX1 \RAM_reg<50><9>  ( .D(\wd<9> ), .E(n18337), .CK(clk), .Q(\RAM<50><9> ) );
  EDFFX1 \RAM_reg<50><8>  ( .D(\wd<8> ), .E(n18337), .CK(clk), .Q(\RAM<50><8> ) );
  EDFFX1 \RAM_reg<50><7>  ( .D(\wd<7> ), .E(n3553), .CK(clk), .Q(\RAM<50><7> )
         );
  EDFFX1 \RAM_reg<50><6>  ( .D(\wd<6> ), .E(n3553), .CK(clk), .Q(\RAM<50><6> )
         );
  EDFFX1 \RAM_reg<50><5>  ( .D(\wd<5> ), .E(n18336), .CK(clk), .Q(\RAM<50><5> ) );
  EDFFX1 \RAM_reg<50><4>  ( .D(\wd<4> ), .E(n18337), .CK(clk), .Q(\RAM<50><4> ) );
  EDFFX1 \RAM_reg<50><3>  ( .D(\wd<3> ), .E(n18336), .CK(clk), .Q(\RAM<50><3> ) );
  EDFFX1 \RAM_reg<50><2>  ( .D(\wd<2> ), .E(n18337), .CK(clk), .Q(\RAM<50><2> ) );
  EDFFX1 \RAM_reg<50><1>  ( .D(\wd<1> ), .E(n18336), .CK(clk), .Q(\RAM<50><1> ) );
  EDFFX1 \RAM_reg<50><0>  ( .D(\wd<0> ), .E(n18337), .CK(clk), .Q(\RAM<50><0> ) );
  EDFFX1 \RAM_reg<42><31>  ( .D(\wd<31> ), .E(n18387), .CK(clk), .Q(
        \RAM<42><31> ) );
  EDFFX1 \RAM_reg<42><30>  ( .D(\wd<30> ), .E(n18387), .CK(clk), .Q(
        \RAM<42><30> ) );
  EDFFX1 \RAM_reg<42><29>  ( .D(\wd<29> ), .E(n18387), .CK(clk), .Q(
        \RAM<42><29> ) );
  EDFFX1 \RAM_reg<42><28>  ( .D(\wd<28> ), .E(n18387), .CK(clk), .Q(
        \RAM<42><28> ) );
  EDFFX1 \RAM_reg<42><27>  ( .D(\wd<27> ), .E(n18387), .CK(clk), .Q(
        \RAM<42><27> ) );
  EDFFX1 \RAM_reg<42><26>  ( .D(\wd<26> ), .E(n18387), .CK(clk), .Q(
        \RAM<42><26> ) );
  EDFFX1 \RAM_reg<42><25>  ( .D(\wd<25> ), .E(n18387), .CK(clk), .Q(
        \RAM<42><25> ) );
  EDFFX1 \RAM_reg<42><24>  ( .D(\wd<24> ), .E(n18387), .CK(clk), .Q(
        \RAM<42><24> ) );
  EDFFX1 \RAM_reg<42><23>  ( .D(\wd<23> ), .E(n18387), .CK(clk), .Q(
        \RAM<42><23> ) );
  EDFFX1 \RAM_reg<42><22>  ( .D(\wd<22> ), .E(n18387), .CK(clk), .Q(
        \RAM<42><22> ) );
  EDFFX1 \RAM_reg<42><21>  ( .D(\wd<21> ), .E(n18387), .CK(clk), .Q(
        \RAM<42><21> ) );
  EDFFX1 \RAM_reg<42><20>  ( .D(\wd<20> ), .E(n18387), .CK(clk), .Q(
        \RAM<42><20> ) );
  EDFFX1 \RAM_reg<42><19>  ( .D(\wd<19> ), .E(n18388), .CK(clk), .Q(
        \RAM<42><19> ) );
  EDFFX1 \RAM_reg<42><18>  ( .D(\wd<18> ), .E(n18388), .CK(clk), .Q(
        \RAM<42><18> ) );
  EDFFX1 \RAM_reg<42><17>  ( .D(\wd<17> ), .E(n18388), .CK(clk), .Q(
        \RAM<42><17> ) );
  EDFFX1 \RAM_reg<42><16>  ( .D(\wd<16> ), .E(n18388), .CK(clk), .Q(
        \RAM<42><16> ) );
  EDFFX1 \RAM_reg<42><15>  ( .D(\wd<15> ), .E(n18388), .CK(clk), .Q(
        \RAM<42><15> ) );
  EDFFX1 \RAM_reg<42><14>  ( .D(\wd<14> ), .E(n18388), .CK(clk), .Q(
        \RAM<42><14> ) );
  EDFFX1 \RAM_reg<42><13>  ( .D(\wd<13> ), .E(n18388), .CK(clk), .Q(
        \RAM<42><13> ) );
  EDFFX1 \RAM_reg<42><12>  ( .D(\wd<12> ), .E(n18388), .CK(clk), .Q(
        \RAM<42><12> ) );
  EDFFX1 \RAM_reg<42><11>  ( .D(\wd<11> ), .E(n18388), .CK(clk), .Q(
        \RAM<42><11> ) );
  EDFFX1 \RAM_reg<42><10>  ( .D(\wd<10> ), .E(n18388), .CK(clk), .Q(
        \RAM<42><10> ) );
  EDFFX1 \RAM_reg<42><9>  ( .D(\wd<9> ), .E(n18388), .CK(clk), .Q(\RAM<42><9> ) );
  EDFFX1 \RAM_reg<42><8>  ( .D(\wd<8> ), .E(n18388), .CK(clk), .Q(\RAM<42><8> ) );
  EDFFX1 \RAM_reg<42><7>  ( .D(\wd<7> ), .E(n3534), .CK(clk), .Q(\RAM<42><7> )
         );
  EDFFX1 \RAM_reg<42><6>  ( .D(\wd<6> ), .E(n3534), .CK(clk), .Q(\RAM<42><6> )
         );
  EDFFX1 \RAM_reg<42><5>  ( .D(\wd<5> ), .E(n18387), .CK(clk), .Q(\RAM<42><5> ) );
  EDFFX1 \RAM_reg<42><4>  ( .D(\wd<4> ), .E(n18388), .CK(clk), .Q(\RAM<42><4> ) );
  EDFFX1 \RAM_reg<42><3>  ( .D(\wd<3> ), .E(n18387), .CK(clk), .Q(\RAM<42><3> ) );
  EDFFX1 \RAM_reg<42><2>  ( .D(\wd<2> ), .E(n18388), .CK(clk), .Q(\RAM<42><2> ) );
  EDFFX1 \RAM_reg<42><1>  ( .D(\wd<1> ), .E(n18387), .CK(clk), .Q(\RAM<42><1> ) );
  EDFFX1 \RAM_reg<42><0>  ( .D(\wd<0> ), .E(n18388), .CK(clk), .Q(\RAM<42><0> ) );
  EDFFX1 \RAM_reg<34><31>  ( .D(\wd<31> ), .E(n18303), .CK(clk), .Q(
        \RAM<34><31> ) );
  EDFFX1 \RAM_reg<34><30>  ( .D(\wd<30> ), .E(n18303), .CK(clk), .Q(
        \RAM<34><30> ) );
  EDFFX1 \RAM_reg<34><29>  ( .D(\wd<29> ), .E(n18303), .CK(clk), .Q(
        \RAM<34><29> ) );
  EDFFX1 \RAM_reg<34><28>  ( .D(\wd<28> ), .E(n18303), .CK(clk), .Q(
        \RAM<34><28> ) );
  EDFFX1 \RAM_reg<34><27>  ( .D(\wd<27> ), .E(n18303), .CK(clk), .Q(
        \RAM<34><27> ) );
  EDFFX1 \RAM_reg<34><26>  ( .D(\wd<26> ), .E(n18303), .CK(clk), .Q(
        \RAM<34><26> ) );
  EDFFX1 \RAM_reg<34><25>  ( .D(\wd<25> ), .E(n18303), .CK(clk), .Q(
        \RAM<34><25> ) );
  EDFFX1 \RAM_reg<34><24>  ( .D(\wd<24> ), .E(n18303), .CK(clk), .Q(
        \RAM<34><24> ) );
  EDFFX1 \RAM_reg<34><23>  ( .D(\wd<23> ), .E(n18303), .CK(clk), .Q(
        \RAM<34><23> ) );
  EDFFX1 \RAM_reg<34><22>  ( .D(\wd<22> ), .E(n18303), .CK(clk), .Q(
        \RAM<34><22> ) );
  EDFFX1 \RAM_reg<34><21>  ( .D(\wd<21> ), .E(n18303), .CK(clk), .Q(
        \RAM<34><21> ) );
  EDFFX1 \RAM_reg<34><20>  ( .D(\wd<20> ), .E(n18303), .CK(clk), .Q(
        \RAM<34><20> ) );
  EDFFX1 \RAM_reg<34><19>  ( .D(\wd<19> ), .E(n18304), .CK(clk), .Q(
        \RAM<34><19> ) );
  EDFFX1 \RAM_reg<34><18>  ( .D(\wd<18> ), .E(n18304), .CK(clk), .Q(
        \RAM<34><18> ) );
  EDFFX1 \RAM_reg<34><17>  ( .D(\wd<17> ), .E(n18304), .CK(clk), .Q(
        \RAM<34><17> ) );
  EDFFX1 \RAM_reg<34><16>  ( .D(\wd<16> ), .E(n18304), .CK(clk), .Q(
        \RAM<34><16> ) );
  EDFFX1 \RAM_reg<34><15>  ( .D(\wd<15> ), .E(n18304), .CK(clk), .Q(
        \RAM<34><15> ) );
  EDFFX1 \RAM_reg<34><14>  ( .D(\wd<14> ), .E(n18304), .CK(clk), .Q(
        \RAM<34><14> ) );
  EDFFX1 \RAM_reg<34><13>  ( .D(\wd<13> ), .E(n18304), .CK(clk), .Q(
        \RAM<34><13> ) );
  EDFFX1 \RAM_reg<34><12>  ( .D(\wd<12> ), .E(n18304), .CK(clk), .Q(
        \RAM<34><12> ) );
  EDFFX1 \RAM_reg<34><11>  ( .D(\wd<11> ), .E(n18304), .CK(clk), .Q(
        \RAM<34><11> ) );
  EDFFX1 \RAM_reg<34><10>  ( .D(\wd<10> ), .E(n18304), .CK(clk), .Q(
        \RAM<34><10> ) );
  EDFFX1 \RAM_reg<34><9>  ( .D(\wd<9> ), .E(n18304), .CK(clk), .Q(\RAM<34><9> ) );
  EDFFX1 \RAM_reg<34><8>  ( .D(\wd<8> ), .E(n18304), .CK(clk), .Q(\RAM<34><8> ) );
  EDFFX1 \RAM_reg<34><7>  ( .D(\wd<7> ), .E(n3568), .CK(clk), .Q(\RAM<34><7> )
         );
  EDFFX1 \RAM_reg<34><6>  ( .D(\wd<6> ), .E(n3568), .CK(clk), .Q(\RAM<34><6> )
         );
  EDFFX1 \RAM_reg<34><5>  ( .D(\wd<5> ), .E(n18303), .CK(clk), .Q(\RAM<34><5> ) );
  EDFFX1 \RAM_reg<34><4>  ( .D(\wd<4> ), .E(n18304), .CK(clk), .Q(\RAM<34><4> ) );
  EDFFX1 \RAM_reg<34><3>  ( .D(\wd<3> ), .E(n18303), .CK(clk), .Q(\RAM<34><3> ) );
  EDFFX1 \RAM_reg<34><2>  ( .D(\wd<2> ), .E(n18304), .CK(clk), .Q(\RAM<34><2> ) );
  EDFFX1 \RAM_reg<34><1>  ( .D(\wd<1> ), .E(n18303), .CK(clk), .Q(\RAM<34><1> ) );
  EDFFX1 \RAM_reg<34><0>  ( .D(\wd<0> ), .E(n18304), .CK(clk), .Q(\RAM<34><0> ) );
  EDFFX1 \RAM_reg<26><31>  ( .D(n18563), .E(n18258), .CK(clk), .Q(
        \RAM<26><31> ) );
  EDFFX1 \RAM_reg<26><30>  ( .D(n18559), .E(n18258), .CK(clk), .Q(
        \RAM<26><30> ) );
  EDFFX1 \RAM_reg<26><29>  ( .D(n18555), .E(n18258), .CK(clk), .Q(
        \RAM<26><29> ) );
  EDFFX1 \RAM_reg<26><28>  ( .D(n18551), .E(n18258), .CK(clk), .Q(
        \RAM<26><28> ) );
  EDFFX1 \RAM_reg<26><27>  ( .D(n18547), .E(n18258), .CK(clk), .Q(
        \RAM<26><27> ) );
  EDFFX1 \RAM_reg<26><26>  ( .D(n18543), .E(n18258), .CK(clk), .Q(
        \RAM<26><26> ) );
  EDFFX1 \RAM_reg<26><25>  ( .D(n18539), .E(n18258), .CK(clk), .Q(
        \RAM<26><25> ) );
  EDFFX1 \RAM_reg<26><24>  ( .D(n18535), .E(n18258), .CK(clk), .Q(
        \RAM<26><24> ) );
  EDFFX1 \RAM_reg<26><23>  ( .D(n18531), .E(n18258), .CK(clk), .Q(
        \RAM<26><23> ) );
  EDFFX1 \RAM_reg<26><22>  ( .D(n18527), .E(n18258), .CK(clk), .Q(
        \RAM<26><22> ) );
  EDFFX1 \RAM_reg<26><21>  ( .D(n18523), .E(n18258), .CK(clk), .Q(
        \RAM<26><21> ) );
  EDFFX1 \RAM_reg<26><20>  ( .D(n18519), .E(n18258), .CK(clk), .Q(
        \RAM<26><20> ) );
  EDFFX1 \RAM_reg<26><19>  ( .D(n18515), .E(n18259), .CK(clk), .Q(
        \RAM<26><19> ) );
  EDFFX1 \RAM_reg<26><18>  ( .D(n18511), .E(n18259), .CK(clk), .Q(
        \RAM<26><18> ) );
  EDFFX1 \RAM_reg<26><17>  ( .D(n18507), .E(n18259), .CK(clk), .Q(
        \RAM<26><17> ) );
  EDFFX1 \RAM_reg<26><16>  ( .D(n18503), .E(n18259), .CK(clk), .Q(
        \RAM<26><16> ) );
  EDFFX1 \RAM_reg<26><15>  ( .D(n18499), .E(n18259), .CK(clk), .Q(
        \RAM<26><15> ) );
  EDFFX1 \RAM_reg<26><14>  ( .D(n18495), .E(n18259), .CK(clk), .Q(
        \RAM<26><14> ) );
  EDFFX1 \RAM_reg<26><13>  ( .D(n18491), .E(n18259), .CK(clk), .Q(
        \RAM<26><13> ) );
  EDFFX1 \RAM_reg<26><12>  ( .D(n18487), .E(n18259), .CK(clk), .Q(
        \RAM<26><12> ) );
  EDFFX1 \RAM_reg<26><11>  ( .D(n18483), .E(n18259), .CK(clk), .Q(
        \RAM<26><11> ) );
  EDFFX1 \RAM_reg<26><10>  ( .D(n18479), .E(n18259), .CK(clk), .Q(
        \RAM<26><10> ) );
  EDFFX1 \RAM_reg<26><9>  ( .D(n18475), .E(n18259), .CK(clk), .Q(\RAM<26><9> )
         );
  EDFFX1 \RAM_reg<26><8>  ( .D(n18471), .E(n18259), .CK(clk), .Q(\RAM<26><8> )
         );
  EDFFX1 \RAM_reg<26><7>  ( .D(n18467), .E(n3583), .CK(clk), .Q(\RAM<26><7> )
         );
  EDFFX1 \RAM_reg<26><6>  ( .D(n18463), .E(n3583), .CK(clk), .Q(\RAM<26><6> )
         );
  EDFFX1 \RAM_reg<26><5>  ( .D(n18459), .E(n18258), .CK(clk), .Q(\RAM<26><5> )
         );
  EDFFX1 \RAM_reg<26><4>  ( .D(n18455), .E(n18259), .CK(clk), .Q(\RAM<26><4> )
         );
  EDFFX1 \RAM_reg<26><3>  ( .D(n18451), .E(n18258), .CK(clk), .Q(\RAM<26><3> )
         );
  EDFFX1 \RAM_reg<26><2>  ( .D(n18447), .E(n18259), .CK(clk), .Q(\RAM<26><2> )
         );
  EDFFX1 \RAM_reg<26><1>  ( .D(n18443), .E(n18258), .CK(clk), .Q(\RAM<26><1> )
         );
  EDFFX1 \RAM_reg<26><0>  ( .D(n18439), .E(n18259), .CK(clk), .Q(\RAM<26><0> )
         );
  EDFFX1 \RAM_reg<18><31>  ( .D(n18564), .E(n18261), .CK(clk), .Q(
        \RAM<18><31> ) );
  EDFFX1 \RAM_reg<18><30>  ( .D(n18560), .E(n18261), .CK(clk), .Q(
        \RAM<18><30> ) );
  EDFFX1 \RAM_reg<18><29>  ( .D(n18556), .E(n18261), .CK(clk), .Q(
        \RAM<18><29> ) );
  EDFFX1 \RAM_reg<18><28>  ( .D(n18552), .E(n18261), .CK(clk), .Q(
        \RAM<18><28> ) );
  EDFFX1 \RAM_reg<18><27>  ( .D(n18548), .E(n18261), .CK(clk), .Q(
        \RAM<18><27> ) );
  EDFFX1 \RAM_reg<18><26>  ( .D(n18544), .E(n18261), .CK(clk), .Q(
        \RAM<18><26> ) );
  EDFFX1 \RAM_reg<18><25>  ( .D(n18540), .E(n18261), .CK(clk), .Q(
        \RAM<18><25> ) );
  EDFFX1 \RAM_reg<18><24>  ( .D(n18536), .E(n18261), .CK(clk), .Q(
        \RAM<18><24> ) );
  EDFFX1 \RAM_reg<18><23>  ( .D(n18532), .E(n18261), .CK(clk), .Q(
        \RAM<18><23> ) );
  EDFFX1 \RAM_reg<18><22>  ( .D(n18528), .E(n18261), .CK(clk), .Q(
        \RAM<18><22> ) );
  EDFFX1 \RAM_reg<18><21>  ( .D(n18524), .E(n18261), .CK(clk), .Q(
        \RAM<18><21> ) );
  EDFFX1 \RAM_reg<18><20>  ( .D(n18520), .E(n18261), .CK(clk), .Q(
        \RAM<18><20> ) );
  EDFFX1 \RAM_reg<18><19>  ( .D(n18516), .E(n18262), .CK(clk), .Q(
        \RAM<18><19> ) );
  EDFFX1 \RAM_reg<18><18>  ( .D(n18512), .E(n18262), .CK(clk), .Q(
        \RAM<18><18> ) );
  EDFFX1 \RAM_reg<18><17>  ( .D(n18508), .E(n18262), .CK(clk), .Q(
        \RAM<18><17> ) );
  EDFFX1 \RAM_reg<18><16>  ( .D(n18504), .E(n18262), .CK(clk), .Q(
        \RAM<18><16> ) );
  EDFFX1 \RAM_reg<18><15>  ( .D(n18500), .E(n18262), .CK(clk), .Q(
        \RAM<18><15> ) );
  EDFFX1 \RAM_reg<18><14>  ( .D(n18496), .E(n18262), .CK(clk), .Q(
        \RAM<18><14> ) );
  EDFFX1 \RAM_reg<18><13>  ( .D(n18492), .E(n18262), .CK(clk), .Q(
        \RAM<18><13> ) );
  EDFFX1 \RAM_reg<18><12>  ( .D(n18488), .E(n18262), .CK(clk), .Q(
        \RAM<18><12> ) );
  EDFFX1 \RAM_reg<18><11>  ( .D(n18484), .E(n18262), .CK(clk), .Q(
        \RAM<18><11> ) );
  EDFFX1 \RAM_reg<18><10>  ( .D(n18480), .E(n18262), .CK(clk), .Q(
        \RAM<18><10> ) );
  EDFFX1 \RAM_reg<18><9>  ( .D(n18476), .E(n18262), .CK(clk), .Q(\RAM<18><9> )
         );
  EDFFX1 \RAM_reg<18><8>  ( .D(n18472), .E(n18262), .CK(clk), .Q(\RAM<18><8> )
         );
  EDFFX1 \RAM_reg<18><7>  ( .D(n18468), .E(n3582), .CK(clk), .Q(\RAM<18><7> )
         );
  EDFFX1 \RAM_reg<18><6>  ( .D(n18464), .E(n3582), .CK(clk), .Q(\RAM<18><6> )
         );
  EDFFX1 \RAM_reg<18><5>  ( .D(n18460), .E(n18261), .CK(clk), .Q(\RAM<18><5> )
         );
  EDFFX1 \RAM_reg<18><4>  ( .D(n18456), .E(n18262), .CK(clk), .Q(\RAM<18><4> )
         );
  EDFFX1 \RAM_reg<18><3>  ( .D(n18452), .E(n18261), .CK(clk), .Q(\RAM<18><3> )
         );
  EDFFX1 \RAM_reg<18><2>  ( .D(n18448), .E(n18262), .CK(clk), .Q(\RAM<18><2> )
         );
  EDFFX1 \RAM_reg<18><1>  ( .D(n18444), .E(n18261), .CK(clk), .Q(\RAM<18><1> )
         );
  EDFFX1 \RAM_reg<18><0>  ( .D(n18440), .E(n18262), .CK(clk), .Q(\RAM<18><0> )
         );
  EDFFX1 \RAM_reg<10><31>  ( .D(n18562), .E(n18264), .CK(clk), .Q(
        \RAM<10><31> ) );
  EDFFX1 \RAM_reg<10><30>  ( .D(n18558), .E(n18264), .CK(clk), .Q(
        \RAM<10><30> ) );
  EDFFX1 \RAM_reg<10><29>  ( .D(n18554), .E(n18264), .CK(clk), .Q(
        \RAM<10><29> ) );
  EDFFX1 \RAM_reg<10><28>  ( .D(n18550), .E(n18264), .CK(clk), .Q(
        \RAM<10><28> ) );
  EDFFX1 \RAM_reg<10><27>  ( .D(n18546), .E(n18264), .CK(clk), .Q(
        \RAM<10><27> ) );
  EDFFX1 \RAM_reg<10><26>  ( .D(n18542), .E(n18264), .CK(clk), .Q(
        \RAM<10><26> ) );
  EDFFX1 \RAM_reg<10><25>  ( .D(n18538), .E(n18264), .CK(clk), .Q(
        \RAM<10><25> ) );
  EDFFX1 \RAM_reg<10><24>  ( .D(n18534), .E(n18264), .CK(clk), .Q(
        \RAM<10><24> ) );
  EDFFX1 \RAM_reg<10><23>  ( .D(n18530), .E(n18264), .CK(clk), .Q(
        \RAM<10><23> ) );
  EDFFX1 \RAM_reg<10><22>  ( .D(n18526), .E(n18264), .CK(clk), .Q(
        \RAM<10><22> ) );
  EDFFX1 \RAM_reg<10><21>  ( .D(n18522), .E(n18264), .CK(clk), .Q(
        \RAM<10><21> ) );
  EDFFX1 \RAM_reg<10><20>  ( .D(n18518), .E(n18264), .CK(clk), .Q(
        \RAM<10><20> ) );
  EDFFX1 \RAM_reg<10><19>  ( .D(n18514), .E(n18265), .CK(clk), .Q(
        \RAM<10><19> ) );
  EDFFX1 \RAM_reg<10><18>  ( .D(n18510), .E(n18265), .CK(clk), .Q(
        \RAM<10><18> ) );
  EDFFX1 \RAM_reg<10><17>  ( .D(n18506), .E(n18265), .CK(clk), .Q(
        \RAM<10><17> ) );
  EDFFX1 \RAM_reg<10><16>  ( .D(n18502), .E(n18265), .CK(clk), .Q(
        \RAM<10><16> ) );
  EDFFX1 \RAM_reg<10><15>  ( .D(n18498), .E(n18265), .CK(clk), .Q(
        \RAM<10><15> ) );
  EDFFX1 \RAM_reg<10><14>  ( .D(n18494), .E(n18265), .CK(clk), .Q(
        \RAM<10><14> ) );
  EDFFX1 \RAM_reg<10><13>  ( .D(n18490), .E(n18265), .CK(clk), .Q(
        \RAM<10><13> ) );
  EDFFX1 \RAM_reg<10><12>  ( .D(n18486), .E(n18265), .CK(clk), .Q(
        \RAM<10><12> ) );
  EDFFX1 \RAM_reg<10><11>  ( .D(n18482), .E(n18265), .CK(clk), .Q(
        \RAM<10><11> ) );
  EDFFX1 \RAM_reg<10><10>  ( .D(n18478), .E(n18265), .CK(clk), .Q(
        \RAM<10><10> ) );
  EDFFX1 \RAM_reg<10><9>  ( .D(n18474), .E(n18265), .CK(clk), .Q(\RAM<10><9> )
         );
  EDFFX1 \RAM_reg<10><8>  ( .D(n18470), .E(n18265), .CK(clk), .Q(\RAM<10><8> )
         );
  EDFFX1 \RAM_reg<10><7>  ( .D(n18466), .E(n3569), .CK(clk), .Q(\RAM<10><7> )
         );
  EDFFX1 \RAM_reg<10><6>  ( .D(n18462), .E(n3569), .CK(clk), .Q(\RAM<10><6> )
         );
  EDFFX1 \RAM_reg<10><5>  ( .D(n18458), .E(n18264), .CK(clk), .Q(\RAM<10><5> )
         );
  EDFFX1 \RAM_reg<10><4>  ( .D(n18454), .E(n18265), .CK(clk), .Q(\RAM<10><4> )
         );
  EDFFX1 \RAM_reg<10><3>  ( .D(n18450), .E(n18264), .CK(clk), .Q(\RAM<10><3> )
         );
  EDFFX1 \RAM_reg<10><2>  ( .D(n18446), .E(n18265), .CK(clk), .Q(\RAM<10><2> )
         );
  EDFFX1 \RAM_reg<10><1>  ( .D(n18442), .E(n18264), .CK(clk), .Q(\RAM<10><1> )
         );
  EDFFX1 \RAM_reg<10><0>  ( .D(n18438), .E(n18265), .CK(clk), .Q(\RAM<10><0> )
         );
  EDFFX1 \RAM_reg<2><31>  ( .D(n18563), .E(n18267), .CK(clk), .Q(\RAM<2><31> )
         );
  EDFFX1 \RAM_reg<2><30>  ( .D(n18559), .E(n18267), .CK(clk), .Q(\RAM<2><30> )
         );
  EDFFX1 \RAM_reg<2><29>  ( .D(n18555), .E(n18267), .CK(clk), .Q(\RAM<2><29> )
         );
  EDFFX1 \RAM_reg<2><28>  ( .D(n18551), .E(n18267), .CK(clk), .Q(\RAM<2><28> )
         );
  EDFFX1 \RAM_reg<2><27>  ( .D(n18547), .E(n18267), .CK(clk), .Q(\RAM<2><27> )
         );
  EDFFX1 \RAM_reg<2><26>  ( .D(n18543), .E(n18267), .CK(clk), .Q(\RAM<2><26> )
         );
  EDFFX1 \RAM_reg<2><25>  ( .D(n18539), .E(n18267), .CK(clk), .Q(\RAM<2><25> )
         );
  EDFFX1 \RAM_reg<2><24>  ( .D(n18535), .E(n18267), .CK(clk), .Q(\RAM<2><24> )
         );
  EDFFX1 \RAM_reg<2><23>  ( .D(n18531), .E(n18267), .CK(clk), .Q(\RAM<2><23> )
         );
  EDFFX1 \RAM_reg<2><22>  ( .D(n18527), .E(n18267), .CK(clk), .Q(\RAM<2><22> )
         );
  EDFFX1 \RAM_reg<2><21>  ( .D(n18523), .E(n18267), .CK(clk), .Q(\RAM<2><21> )
         );
  EDFFX1 \RAM_reg<2><20>  ( .D(n18519), .E(n18267), .CK(clk), .Q(\RAM<2><20> )
         );
  EDFFX1 \RAM_reg<2><19>  ( .D(n18515), .E(n18268), .CK(clk), .Q(\RAM<2><19> )
         );
  EDFFX1 \RAM_reg<2><18>  ( .D(n18511), .E(n18268), .CK(clk), .Q(\RAM<2><18> )
         );
  EDFFX1 \RAM_reg<2><17>  ( .D(n18507), .E(n18268), .CK(clk), .Q(\RAM<2><17> )
         );
  EDFFX1 \RAM_reg<2><16>  ( .D(n18503), .E(n18268), .CK(clk), .Q(\RAM<2><16> )
         );
  EDFFX1 \RAM_reg<2><15>  ( .D(n18499), .E(n18268), .CK(clk), .Q(\RAM<2><15> )
         );
  EDFFX1 \RAM_reg<2><14>  ( .D(n18495), .E(n18268), .CK(clk), .Q(\RAM<2><14> )
         );
  EDFFX1 \RAM_reg<2><13>  ( .D(n18491), .E(n18268), .CK(clk), .Q(\RAM<2><13> )
         );
  EDFFX1 \RAM_reg<2><12>  ( .D(n18487), .E(n18268), .CK(clk), .Q(\RAM<2><12> )
         );
  EDFFX1 \RAM_reg<2><11>  ( .D(n18483), .E(n18268), .CK(clk), .Q(\RAM<2><11> )
         );
  EDFFX1 \RAM_reg<2><10>  ( .D(n18479), .E(n18268), .CK(clk), .Q(\RAM<2><10> )
         );
  EDFFX1 \RAM_reg<2><9>  ( .D(n18475), .E(n18268), .CK(clk), .Q(\RAM<2><9> )
         );
  EDFFX1 \RAM_reg<2><8>  ( .D(n18471), .E(n18268), .CK(clk), .Q(\RAM<2><8> )
         );
  EDFFX1 \RAM_reg<2><7>  ( .D(n18467), .E(n3565), .CK(clk), .Q(\RAM<2><7> ) );
  EDFFX1 \RAM_reg<2><6>  ( .D(n18463), .E(n3565), .CK(clk), .Q(\RAM<2><6> ) );
  EDFFX1 \RAM_reg<2><5>  ( .D(n18459), .E(n18267), .CK(clk), .Q(\RAM<2><5> )
         );
  EDFFX1 \RAM_reg<2><4>  ( .D(n18455), .E(n18268), .CK(clk), .Q(\RAM<2><4> )
         );
  EDFFX1 \RAM_reg<2><3>  ( .D(n18451), .E(n18267), .CK(clk), .Q(\RAM<2><3> )
         );
  EDFFX1 \RAM_reg<2><2>  ( .D(n18447), .E(n18268), .CK(clk), .Q(\RAM<2><2> )
         );
  EDFFX1 \RAM_reg<2><1>  ( .D(n18443), .E(n18267), .CK(clk), .Q(\RAM<2><1> )
         );
  EDFFX1 \RAM_reg<2><0>  ( .D(n18439), .E(n18268), .CK(clk), .Q(\RAM<2><0> )
         );
  OR2X2 U2 ( .A(n18566), .B(N36), .Y(n16074) );
  OR2X2 U3 ( .A(n18566), .B(n18567), .Y(n16075) );
  OR2X2 U4 ( .A(n18567), .B(N37), .Y(n16076) );
  OR2X2 U5 ( .A(N37), .B(N36), .Y(n16077) );
  CLKINVX3 U6 ( .A(n18257), .Y(n18256) );
  CLKINVX3 U7 ( .A(n18254), .Y(n18253) );
  CLKINVX3 U8 ( .A(n18251), .Y(n18250) );
  CLKINVX3 U9 ( .A(n18248), .Y(n18247) );
  CLKINVX3 U10 ( .A(n18413), .Y(n18412) );
  CLKINVX3 U11 ( .A(n18419), .Y(n18418) );
  CLKINVX3 U12 ( .A(n18350), .Y(n18349) );
  CLKINVX3 U13 ( .A(n18359), .Y(n18358) );
  CLKINVX3 U14 ( .A(n18335), .Y(n18334) );
  CLKINVX3 U15 ( .A(n18278), .Y(n18277) );
  CLKINVX3 U16 ( .A(n18308), .Y(n18307) );
  CLKINVX3 U17 ( .A(n18275), .Y(n18274) );
  CLKINVX3 U18 ( .A(n18311), .Y(n18310) );
  CLKINVX3 U19 ( .A(n18434), .Y(n18433) );
  CLKINVX3 U20 ( .A(n18431), .Y(n18430) );
  CLKINVX3 U21 ( .A(n18368), .Y(n18367) );
  CLKINVX3 U22 ( .A(n18395), .Y(n18394) );
  CLKINVX3 U23 ( .A(n18317), .Y(n18316) );
  CLKINVX3 U24 ( .A(n18398), .Y(n18397) );
  CLKINVX3 U25 ( .A(n18281), .Y(n18280) );
  CLKINVX3 U26 ( .A(n18383), .Y(n18382) );
  CLKINVX3 U27 ( .A(n18344), .Y(n18343) );
  CLKINVX3 U28 ( .A(n18326), .Y(n18325) );
  CLKINVX3 U29 ( .A(n18272), .Y(n18271) );
  CLKINVX3 U30 ( .A(n18299), .Y(n18298) );
  CLKINVX3 U31 ( .A(n18293), .Y(n18292) );
  CLKINVX3 U32 ( .A(n18374), .Y(n18373) );
  CLKINVX3 U33 ( .A(n18428), .Y(n18427) );
  CLKINVX3 U34 ( .A(n18341), .Y(n18340) );
  CLKINVX3 U35 ( .A(n18386), .Y(n18385) );
  CLKINVX3 U36 ( .A(n18392), .Y(n18391) );
  CLKINVX3 U37 ( .A(n18329), .Y(n18328) );
  CLKINVX3 U38 ( .A(n18269), .Y(n18268) );
  CLKINVX3 U39 ( .A(n18266), .Y(n18265) );
  CLKINVX3 U40 ( .A(n18263), .Y(n18262) );
  CLKINVX3 U41 ( .A(n18260), .Y(n18259) );
  CLKINVX3 U42 ( .A(n18305), .Y(n18304) );
  CLKINVX3 U43 ( .A(n18389), .Y(n18388) );
  CLKINVX3 U44 ( .A(n18338), .Y(n18337) );
  CLKINVX3 U45 ( .A(n18332), .Y(n18331) );
  CLKINVX3 U46 ( .A(n18290), .Y(n18289) );
  CLKINVX3 U47 ( .A(n18437), .Y(n18436) );
  CLKINVX3 U48 ( .A(n18284), .Y(n18283) );
  CLKINVX3 U49 ( .A(n18320), .Y(n18319) );
  CLKINVX3 U50 ( .A(n18425), .Y(n18424) );
  CLKINVX3 U51 ( .A(n18314), .Y(n18313) );
  CLKINVX3 U52 ( .A(n18422), .Y(n18421) );
  CLKINVX3 U53 ( .A(n18380), .Y(n18379) );
  CLKINVX3 U54 ( .A(n18401), .Y(n18400) );
  CLKINVX3 U55 ( .A(n18410), .Y(n18409) );
  CLKINVX3 U56 ( .A(n18404), .Y(n18403) );
  CLKINVX3 U57 ( .A(n18407), .Y(n18406) );
  CLKINVX3 U58 ( .A(n18323), .Y(n18322) );
  CLKINVX3 U59 ( .A(n18353), .Y(n18352) );
  CLKINVX3 U60 ( .A(n18362), .Y(n18361) );
  CLKINVX3 U61 ( .A(n18356), .Y(n18355) );
  CLKINVX3 U62 ( .A(n18302), .Y(n18301) );
  CLKINVX3 U63 ( .A(n18287), .Y(n18286) );
  CLKINVX3 U64 ( .A(n18371), .Y(n18370) );
  CLKINVX3 U65 ( .A(n18296), .Y(n18295) );
  CLKINVX3 U66 ( .A(n18416), .Y(n18415) );
  CLKINVX3 U67 ( .A(n18377), .Y(n18376) );
  CLKINVX3 U68 ( .A(n18347), .Y(n18346) );
  CLKINVX3 U69 ( .A(n18365), .Y(n18364) );
  CLKINVX3 U70 ( .A(n18145), .Y(n18144) );
  CLKINVX3 U71 ( .A(n18145), .Y(n18140) );
  CLKINVX3 U72 ( .A(n18145), .Y(n18141) );
  CLKINVX3 U73 ( .A(n18145), .Y(n18142) );
  CLKINVX3 U74 ( .A(n18145), .Y(n18143) );
  CLKINVX3 U75 ( .A(n18275), .Y(n18273) );
  INVX1 U76 ( .A(n3580), .Y(n18275) );
  CLKINVX3 U77 ( .A(n18269), .Y(n18267) );
  INVX1 U78 ( .A(n3565), .Y(n18269) );
  CLKINVX3 U79 ( .A(n18257), .Y(n18255) );
  INVX1 U80 ( .A(n3560), .Y(n18257) );
  CLKINVX3 U81 ( .A(n18434), .Y(n18432) );
  INVX1 U82 ( .A(n3519), .Y(n18434) );
  CLKINVX3 U83 ( .A(n18368), .Y(n18366) );
  INVX1 U84 ( .A(n3542), .Y(n18368) );
  CLKINVX3 U85 ( .A(n18281), .Y(n18279) );
  INVX1 U86 ( .A(n3578), .Y(n18281) );
  CLKINVX3 U87 ( .A(n18272), .Y(n18270) );
  INVX1 U88 ( .A(n3581), .Y(n18272) );
  CLKINVX3 U89 ( .A(n18266), .Y(n18264) );
  INVX1 U90 ( .A(n3569), .Y(n18266) );
  CLKINVX3 U91 ( .A(n18263), .Y(n18261) );
  INVX1 U92 ( .A(n3582), .Y(n18263) );
  CLKINVX3 U93 ( .A(n18260), .Y(n18258) );
  INVX1 U94 ( .A(n3583), .Y(n18260) );
  CLKINVX3 U95 ( .A(n18389), .Y(n18387) );
  INVX1 U96 ( .A(n3534), .Y(n18389) );
  CLKINVX3 U97 ( .A(n18332), .Y(n18330) );
  INVX1 U98 ( .A(n3555), .Y(n18332) );
  CLKINVX3 U99 ( .A(n18437), .Y(n18435) );
  INVX1 U100 ( .A(n66), .Y(n18437) );
  CLKINVX3 U101 ( .A(n18320), .Y(n18318) );
  INVX1 U102 ( .A(n3559), .Y(n18320) );
  CLKINVX3 U103 ( .A(n18314), .Y(n18312) );
  INVX1 U104 ( .A(n3563), .Y(n18314) );
  CLKINVX3 U105 ( .A(n18380), .Y(n18378) );
  INVX1 U106 ( .A(n3538), .Y(n18380) );
  CLKINVX3 U107 ( .A(n18407), .Y(n18405) );
  INVX1 U108 ( .A(n3528), .Y(n18407) );
  CLKINVX3 U109 ( .A(n18356), .Y(n18354) );
  INVX1 U110 ( .A(n3546), .Y(n18356) );
  CLKINVX3 U111 ( .A(n18254), .Y(n18252) );
  INVX1 U112 ( .A(n3561), .Y(n18254) );
  CLKINVX3 U113 ( .A(n18251), .Y(n18249) );
  INVX1 U114 ( .A(n3566), .Y(n18251) );
  CLKINVX3 U115 ( .A(n18248), .Y(n18246) );
  INVX1 U116 ( .A(n3576), .Y(n18248) );
  CLKINVX3 U117 ( .A(n18278), .Y(n18276) );
  INVX1 U118 ( .A(n3579), .Y(n18278) );
  CLKINVX3 U119 ( .A(n18413), .Y(n18411) );
  INVX1 U120 ( .A(n3526), .Y(n18413) );
  CLKINVX3 U121 ( .A(n18419), .Y(n18417) );
  INVX1 U122 ( .A(n3524), .Y(n18419) );
  CLKINVX3 U123 ( .A(n18350), .Y(n18348) );
  INVX1 U124 ( .A(n3549), .Y(n18350) );
  CLKINVX3 U125 ( .A(n18359), .Y(n18357) );
  INVX1 U126 ( .A(n3545), .Y(n18359) );
  CLKINVX3 U127 ( .A(n18335), .Y(n18333) );
  INVX1 U128 ( .A(n3554), .Y(n18335) );
  CLKINVX3 U129 ( .A(n18308), .Y(n18306) );
  INVX1 U130 ( .A(n3567), .Y(n18308) );
  CLKINVX3 U131 ( .A(n18311), .Y(n18309) );
  INVX1 U132 ( .A(n3564), .Y(n18311) );
  CLKINVX3 U133 ( .A(n18431), .Y(n18429) );
  INVX1 U134 ( .A(n3520), .Y(n18431) );
  CLKINVX3 U135 ( .A(n18395), .Y(n18393) );
  INVX1 U136 ( .A(n3532), .Y(n18395) );
  CLKINVX3 U137 ( .A(n18317), .Y(n18315) );
  INVX1 U138 ( .A(n3562), .Y(n18317) );
  CLKINVX3 U139 ( .A(n18398), .Y(n18396) );
  INVX1 U140 ( .A(n3531), .Y(n18398) );
  CLKINVX3 U141 ( .A(n18383), .Y(n18381) );
  INVX1 U142 ( .A(n3536), .Y(n18383) );
  CLKINVX3 U143 ( .A(n18344), .Y(n18342) );
  INVX1 U144 ( .A(n3551), .Y(n18344) );
  CLKINVX3 U145 ( .A(n18326), .Y(n18324) );
  INVX1 U146 ( .A(n3557), .Y(n18326) );
  CLKINVX3 U147 ( .A(n18299), .Y(n18297) );
  INVX1 U148 ( .A(n3571), .Y(n18299) );
  CLKINVX3 U149 ( .A(n18293), .Y(n18291) );
  INVX1 U150 ( .A(n3573), .Y(n18293) );
  CLKINVX3 U151 ( .A(n18374), .Y(n18372) );
  INVX1 U152 ( .A(n3540), .Y(n18374) );
  CLKINVX3 U153 ( .A(n18428), .Y(n18426) );
  INVX1 U154 ( .A(n3521), .Y(n18428) );
  CLKINVX3 U155 ( .A(n18341), .Y(n18339) );
  INVX1 U156 ( .A(n3552), .Y(n18341) );
  CLKINVX3 U157 ( .A(n18386), .Y(n18384) );
  INVX1 U158 ( .A(n3535), .Y(n18386) );
  CLKINVX3 U159 ( .A(n18392), .Y(n18390) );
  INVX1 U160 ( .A(n3533), .Y(n18392) );
  CLKINVX3 U161 ( .A(n18329), .Y(n18327) );
  INVX1 U162 ( .A(n3556), .Y(n18329) );
  CLKINVX3 U163 ( .A(n18305), .Y(n18303) );
  INVX1 U164 ( .A(n3568), .Y(n18305) );
  CLKINVX3 U165 ( .A(n18338), .Y(n18336) );
  INVX1 U166 ( .A(n3553), .Y(n18338) );
  CLKINVX3 U167 ( .A(n18290), .Y(n18288) );
  INVX1 U168 ( .A(n3574), .Y(n18290) );
  CLKINVX3 U169 ( .A(n18284), .Y(n18282) );
  INVX1 U170 ( .A(n3577), .Y(n18284) );
  CLKINVX3 U171 ( .A(n18425), .Y(n18423) );
  INVX1 U172 ( .A(n3522), .Y(n18425) );
  CLKINVX3 U173 ( .A(n18422), .Y(n18420) );
  INVX1 U174 ( .A(n3523), .Y(n18422) );
  CLKINVX3 U175 ( .A(n18401), .Y(n18399) );
  INVX1 U176 ( .A(n3530), .Y(n18401) );
  CLKINVX3 U177 ( .A(n18410), .Y(n18408) );
  INVX1 U178 ( .A(n3527), .Y(n18410) );
  CLKINVX3 U179 ( .A(n18404), .Y(n18402) );
  INVX1 U180 ( .A(n3529), .Y(n18404) );
  CLKINVX3 U181 ( .A(n18323), .Y(n18321) );
  INVX1 U182 ( .A(n3558), .Y(n18323) );
  CLKINVX3 U183 ( .A(n18353), .Y(n18351) );
  INVX1 U184 ( .A(n3548), .Y(n18353) );
  CLKINVX3 U185 ( .A(n18362), .Y(n18360) );
  INVX1 U186 ( .A(n3544), .Y(n18362) );
  CLKINVX3 U187 ( .A(n18302), .Y(n18300) );
  INVX1 U188 ( .A(n3570), .Y(n18302) );
  CLKINVX3 U189 ( .A(n18287), .Y(n18285) );
  INVX1 U190 ( .A(n3575), .Y(n18287) );
  CLKINVX3 U191 ( .A(n18371), .Y(n18369) );
  INVX1 U192 ( .A(n3541), .Y(n18371) );
  CLKINVX3 U193 ( .A(n18296), .Y(n18294) );
  INVX1 U194 ( .A(n3572), .Y(n18296) );
  CLKINVX3 U195 ( .A(n18416), .Y(n18414) );
  INVX1 U196 ( .A(n3525), .Y(n18416) );
  CLKINVX3 U197 ( .A(n18377), .Y(n18375) );
  INVX1 U198 ( .A(n3539), .Y(n18377) );
  CLKINVX3 U199 ( .A(n18347), .Y(n18345) );
  INVX1 U200 ( .A(n3550), .Y(n18347) );
  CLKINVX3 U201 ( .A(n18365), .Y(n18363) );
  INVX1 U202 ( .A(n3543), .Y(n18365) );
  CLKINVX3 U203 ( .A(n16075), .Y(n18131) );
  CLKINVX3 U204 ( .A(n18187), .Y(n18186) );
  CLKINVX3 U205 ( .A(n18173), .Y(n18172) );
  CLKINVX3 U206 ( .A(n18159), .Y(n18158) );
  CLKINVX3 U207 ( .A(n18243), .Y(n18242) );
  CLKINVX3 U208 ( .A(n18229), .Y(n18228) );
  CLKINVX3 U209 ( .A(n18201), .Y(n18200) );
  CLKINVX3 U210 ( .A(n18187), .Y(n18181) );
  CLKINVX3 U211 ( .A(n18173), .Y(n18168) );
  CLKINVX3 U212 ( .A(n18159), .Y(n18154) );
  CLKINVX3 U213 ( .A(n18243), .Y(n18237) );
  CLKINVX3 U214 ( .A(n18215), .Y(n18210) );
  CLKINVX3 U215 ( .A(n18229), .Y(n18223) );
  CLKINVX3 U216 ( .A(n18201), .Y(n18195) );
  CLKINVX3 U217 ( .A(n18187), .Y(n18182) );
  CLKINVX3 U218 ( .A(n18173), .Y(n18169) );
  CLKINVX3 U219 ( .A(n18159), .Y(n18155) );
  CLKINVX3 U220 ( .A(n18215), .Y(n18211) );
  CLKINVX3 U221 ( .A(n18229), .Y(n18224) );
  CLKINVX3 U222 ( .A(n18201), .Y(n18196) );
  CLKINVX3 U223 ( .A(n18187), .Y(n18183) );
  CLKINVX3 U224 ( .A(n18173), .Y(n18171) );
  CLKINVX3 U225 ( .A(n18159), .Y(n18157) );
  CLKINVX3 U226 ( .A(n18243), .Y(n18239) );
  CLKINVX3 U227 ( .A(n18215), .Y(n18212) );
  CLKINVX3 U228 ( .A(n18229), .Y(n18225) );
  CLKINVX3 U229 ( .A(n18201), .Y(n18197) );
  CLKINVX3 U230 ( .A(n18215), .Y(n18213) );
  CLKINVX3 U231 ( .A(n18229), .Y(n18226) );
  CLKINVX3 U232 ( .A(n18201), .Y(n18198) );
  CLKINVX3 U233 ( .A(n18187), .Y(n18184) );
  CLKINVX3 U234 ( .A(n18243), .Y(n18240) );
  CLKINVX3 U235 ( .A(n18215), .Y(n18214) );
  CLKINVX3 U236 ( .A(n18229), .Y(n18227) );
  CLKINVX3 U237 ( .A(n18201), .Y(n18199) );
  CLKINVX3 U238 ( .A(n18187), .Y(n18185) );
  CLKINVX3 U239 ( .A(n18243), .Y(n18241) );
  CLKINVX3 U240 ( .A(n18173), .Y(n18170) );
  CLKINVX3 U241 ( .A(n18159), .Y(n18156) );
  CLKINVX3 U242 ( .A(n18243), .Y(n18238) );
  CLKINVX3 U243 ( .A(n18145), .Y(n18139) );
  INVX1 U244 ( .A(n2085), .Y(n18145) );
  CLKINVX3 U245 ( .A(n18180), .Y(n18179) );
  CLKINVX3 U246 ( .A(n18166), .Y(n18165) );
  CLKINVX3 U247 ( .A(n18152), .Y(n18151) );
  CLKINVX3 U248 ( .A(n18138), .Y(n18137) );
  CLKINVX3 U249 ( .A(n18236), .Y(n18235) );
  CLKINVX3 U250 ( .A(n18208), .Y(n18207) );
  CLKINVX3 U251 ( .A(n18222), .Y(n18221) );
  CLKINVX3 U252 ( .A(n18194), .Y(n18193) );
  CLKINVX3 U253 ( .A(n18180), .Y(n18174) );
  CLKINVX3 U254 ( .A(n18166), .Y(n18160) );
  CLKINVX3 U255 ( .A(n18152), .Y(n18146) );
  CLKINVX3 U256 ( .A(n18138), .Y(n18132) );
  CLKINVX3 U257 ( .A(n18236), .Y(n18230) );
  CLKINVX3 U258 ( .A(n18208), .Y(n18202) );
  CLKINVX3 U259 ( .A(n18222), .Y(n18216) );
  CLKINVX3 U260 ( .A(n18194), .Y(n18189) );
  CLKINVX3 U261 ( .A(n18180), .Y(n18175) );
  CLKINVX3 U262 ( .A(n18166), .Y(n18161) );
  CLKINVX3 U263 ( .A(n18152), .Y(n18147) );
  CLKINVX3 U264 ( .A(n18138), .Y(n18133) );
  CLKINVX3 U265 ( .A(n18236), .Y(n18231) );
  CLKINVX3 U266 ( .A(n18208), .Y(n18203) );
  CLKINVX3 U267 ( .A(n18222), .Y(n18217) );
  CLKINVX3 U268 ( .A(n18194), .Y(n18190) );
  CLKINVX3 U269 ( .A(n18180), .Y(n18176) );
  CLKINVX3 U270 ( .A(n18166), .Y(n18162) );
  CLKINVX3 U271 ( .A(n18152), .Y(n18148) );
  CLKINVX3 U272 ( .A(n18138), .Y(n18134) );
  CLKINVX3 U273 ( .A(n18236), .Y(n18232) );
  CLKINVX3 U274 ( .A(n18208), .Y(n18204) );
  CLKINVX3 U275 ( .A(n18222), .Y(n18218) );
  CLKINVX3 U276 ( .A(n18180), .Y(n18177) );
  CLKINVX3 U277 ( .A(n18166), .Y(n18163) );
  CLKINVX3 U278 ( .A(n18152), .Y(n18149) );
  CLKINVX3 U279 ( .A(n18138), .Y(n18135) );
  CLKINVX3 U280 ( .A(n18236), .Y(n18233) );
  CLKINVX3 U281 ( .A(n18208), .Y(n18205) );
  CLKINVX3 U282 ( .A(n18222), .Y(n18219) );
  CLKINVX3 U283 ( .A(n18194), .Y(n18191) );
  CLKINVX3 U284 ( .A(n18166), .Y(n18164) );
  CLKINVX3 U285 ( .A(n18152), .Y(n18150) );
  CLKINVX3 U286 ( .A(n18138), .Y(n18136) );
  CLKINVX3 U287 ( .A(n18236), .Y(n18234) );
  CLKINVX3 U288 ( .A(n18208), .Y(n18206) );
  CLKINVX3 U289 ( .A(n18222), .Y(n18220) );
  CLKINVX3 U290 ( .A(n18180), .Y(n18178) );
  CLKINVX3 U291 ( .A(n18194), .Y(n18192) );
  CLKINVX3 U292 ( .A(n18441), .Y(n18440) );
  CLKINVX3 U293 ( .A(n18445), .Y(n18444) );
  CLKINVX3 U294 ( .A(n18449), .Y(n18448) );
  CLKINVX3 U295 ( .A(n18453), .Y(n18452) );
  CLKINVX3 U296 ( .A(n18457), .Y(n18456) );
  CLKINVX3 U297 ( .A(n18461), .Y(n18460) );
  CLKINVX3 U298 ( .A(n18465), .Y(n18464) );
  CLKINVX3 U299 ( .A(n18469), .Y(n18468) );
  CLKINVX3 U300 ( .A(n18473), .Y(n18472) );
  CLKINVX3 U301 ( .A(n18477), .Y(n18476) );
  CLKINVX3 U302 ( .A(n18481), .Y(n18480) );
  CLKINVX3 U303 ( .A(n18485), .Y(n18484) );
  CLKINVX3 U304 ( .A(n18489), .Y(n18488) );
  CLKINVX3 U305 ( .A(n18493), .Y(n18492) );
  CLKINVX3 U306 ( .A(n18497), .Y(n18496) );
  CLKINVX3 U307 ( .A(n18501), .Y(n18500) );
  CLKINVX3 U308 ( .A(n18505), .Y(n18504) );
  CLKINVX3 U309 ( .A(n18509), .Y(n18508) );
  CLKINVX3 U310 ( .A(n18513), .Y(n18512) );
  CLKINVX3 U311 ( .A(n18517), .Y(n18516) );
  CLKINVX3 U312 ( .A(n18521), .Y(n18520) );
  CLKINVX3 U313 ( .A(n18525), .Y(n18524) );
  CLKINVX3 U314 ( .A(n18529), .Y(n18528) );
  CLKINVX3 U315 ( .A(n18533), .Y(n18532) );
  CLKINVX3 U316 ( .A(n18537), .Y(n18536) );
  CLKINVX3 U317 ( .A(n18541), .Y(n18540) );
  CLKINVX3 U318 ( .A(n18545), .Y(n18544) );
  CLKINVX3 U319 ( .A(n18549), .Y(n18548) );
  CLKINVX3 U320 ( .A(n18553), .Y(n18552) );
  CLKINVX3 U321 ( .A(n18557), .Y(n18556) );
  CLKINVX3 U322 ( .A(n18561), .Y(n18560) );
  CLKINVX3 U323 ( .A(n18565), .Y(n18564) );
  CLKINVX3 U324 ( .A(n18441), .Y(n18439) );
  CLKINVX3 U325 ( .A(n18445), .Y(n18443) );
  CLKINVX3 U326 ( .A(n18449), .Y(n18447) );
  CLKINVX3 U327 ( .A(n18453), .Y(n18451) );
  CLKINVX3 U328 ( .A(n18457), .Y(n18455) );
  CLKINVX3 U329 ( .A(n18461), .Y(n18459) );
  CLKINVX3 U330 ( .A(n18465), .Y(n18463) );
  CLKINVX3 U331 ( .A(n18469), .Y(n18467) );
  CLKINVX3 U332 ( .A(n18473), .Y(n18471) );
  CLKINVX3 U333 ( .A(n18477), .Y(n18475) );
  CLKINVX3 U334 ( .A(n18481), .Y(n18479) );
  CLKINVX3 U335 ( .A(n18485), .Y(n18483) );
  CLKINVX3 U336 ( .A(n18489), .Y(n18487) );
  CLKINVX3 U337 ( .A(n18493), .Y(n18491) );
  CLKINVX3 U338 ( .A(n18497), .Y(n18495) );
  CLKINVX3 U339 ( .A(n18501), .Y(n18499) );
  CLKINVX3 U340 ( .A(n18505), .Y(n18503) );
  CLKINVX3 U341 ( .A(n18509), .Y(n18507) );
  CLKINVX3 U342 ( .A(n18513), .Y(n18511) );
  CLKINVX3 U343 ( .A(n18517), .Y(n18515) );
  CLKINVX3 U344 ( .A(n18521), .Y(n18519) );
  CLKINVX3 U345 ( .A(n18525), .Y(n18523) );
  CLKINVX3 U346 ( .A(n18529), .Y(n18527) );
  CLKINVX3 U347 ( .A(n18533), .Y(n18531) );
  CLKINVX3 U348 ( .A(n18537), .Y(n18535) );
  CLKINVX3 U349 ( .A(n18541), .Y(n18539) );
  CLKINVX3 U350 ( .A(n18545), .Y(n18543) );
  CLKINVX3 U351 ( .A(n18549), .Y(n18547) );
  CLKINVX3 U352 ( .A(n18553), .Y(n18551) );
  CLKINVX3 U353 ( .A(n18557), .Y(n18555) );
  CLKINVX3 U354 ( .A(n18561), .Y(n18559) );
  CLKINVX3 U355 ( .A(n18565), .Y(n18563) );
  CLKINVX3 U356 ( .A(n18441), .Y(n18438) );
  CLKINVX3 U357 ( .A(n18445), .Y(n18442) );
  CLKINVX3 U358 ( .A(n18449), .Y(n18446) );
  CLKINVX3 U359 ( .A(n18453), .Y(n18450) );
  CLKINVX3 U360 ( .A(n18457), .Y(n18454) );
  CLKINVX3 U361 ( .A(n18461), .Y(n18458) );
  CLKINVX3 U362 ( .A(n18465), .Y(n18462) );
  CLKINVX3 U363 ( .A(n18469), .Y(n18466) );
  CLKINVX3 U364 ( .A(n18473), .Y(n18470) );
  CLKINVX3 U365 ( .A(n18477), .Y(n18474) );
  CLKINVX3 U366 ( .A(n18481), .Y(n18478) );
  CLKINVX3 U367 ( .A(n18485), .Y(n18482) );
  CLKINVX3 U368 ( .A(n18489), .Y(n18486) );
  CLKINVX3 U369 ( .A(n18493), .Y(n18490) );
  CLKINVX3 U370 ( .A(n18497), .Y(n18494) );
  CLKINVX3 U371 ( .A(n18501), .Y(n18498) );
  CLKINVX3 U372 ( .A(n18505), .Y(n18502) );
  CLKINVX3 U373 ( .A(n18509), .Y(n18506) );
  CLKINVX3 U374 ( .A(n18513), .Y(n18510) );
  CLKINVX3 U375 ( .A(n18517), .Y(n18514) );
  CLKINVX3 U376 ( .A(n18521), .Y(n18518) );
  CLKINVX3 U377 ( .A(n18525), .Y(n18522) );
  CLKINVX3 U378 ( .A(n18529), .Y(n18526) );
  CLKINVX3 U379 ( .A(n18533), .Y(n18530) );
  CLKINVX3 U380 ( .A(n18537), .Y(n18534) );
  CLKINVX3 U381 ( .A(n18541), .Y(n18538) );
  CLKINVX3 U382 ( .A(n18545), .Y(n18542) );
  CLKINVX3 U383 ( .A(n18549), .Y(n18546) );
  CLKINVX3 U384 ( .A(n18553), .Y(n18550) );
  CLKINVX3 U385 ( .A(n18557), .Y(n18554) );
  CLKINVX3 U386 ( .A(n18561), .Y(n18558) );
  CLKINVX3 U387 ( .A(n18565), .Y(n18562) );
  NAND2X2 U388 ( .A(n3509), .B(n18244), .Y(n3492) );
  NAND2X2 U389 ( .A(n3509), .B(n18126), .Y(n3496) );
  NAND2X2 U390 ( .A(n3509), .B(n18128), .Y(n3505) );
  NAND2X2 U391 ( .A(n3509), .B(n18130), .Y(n3508) );
  NOR2X1 U392 ( .A(n3494), .B(n3499), .Y(n3569) );
  NOR2X1 U393 ( .A(n3494), .B(n3496), .Y(n3582) );
  NOR2X1 U394 ( .A(n3494), .B(n3495), .Y(n3583) );
  NOR2X1 U395 ( .A(n3494), .B(n3505), .Y(n3568) );
  NOR2X1 U396 ( .A(n3494), .B(n3500), .Y(n3534) );
  NOR2X1 U397 ( .A(n3494), .B(n3508), .Y(n3553) );
  NOR2X1 U398 ( .A(n3494), .B(n3497), .Y(n3555) );
  NOR2X1 U399 ( .A(n3493), .B(n3499), .Y(n3559) );
  NOR2X1 U400 ( .A(n3493), .B(n3496), .Y(n3563) );
  NOR2X1 U401 ( .A(n3493), .B(n3495), .Y(n3538) );
  NOR2X1 U402 ( .A(n3493), .B(n3505), .Y(n3527) );
  NOR2X1 U403 ( .A(n3493), .B(n3500), .Y(n3528) );
  NOR2X1 U404 ( .A(n3493), .B(n3508), .Y(n3548) );
  NOR2X1 U405 ( .A(n3493), .B(n3497), .Y(n3546) );
  NOR2X1 U406 ( .A(n3498), .B(n3499), .Y(n3580) );
  NOR2X1 U407 ( .A(n3498), .B(n3505), .Y(n3562) );
  NOR2X1 U408 ( .A(n3498), .B(n3500), .Y(n3578) );
  NOR2X1 U409 ( .A(n3498), .B(n3508), .Y(n3551) );
  NOR2X1 U410 ( .A(n3502), .B(n3505), .Y(n3526) );
  NOR2X1 U411 ( .A(n3502), .B(n3508), .Y(n3549) );
  NOR2X1 U412 ( .A(n3504), .B(n3505), .Y(n3552) );
  NOR2X1 U413 ( .A(n3504), .B(n3508), .Y(n3533) );
  NOR2X1 U414 ( .A(n3501), .B(n3505), .Y(n3530) );
  NOR2X1 U415 ( .A(n3501), .B(n3508), .Y(n3558) );
  NOR2X1 U416 ( .A(n3503), .B(n3505), .Y(n3525) );
  NOR2X1 U417 ( .A(n3503), .B(n3508), .Y(n3550) );
  NOR2X1 U418 ( .A(n3506), .B(n3508), .Y(n3536) );
  NOR2X1 U419 ( .A(n3492), .B(n3502), .Y(n3560) );
  NOR2X1 U420 ( .A(n3492), .B(n3506), .Y(n3554) );
  NOR2X1 U421 ( .A(n3492), .B(n3498), .Y(n3579) );
  NOR2X1 U422 ( .A(n3492), .B(n3504), .Y(n3571) );
  NOR2X1 U423 ( .A(n3492), .B(n3494), .Y(n3565) );
  NOR2X1 U424 ( .A(n3492), .B(n3501), .Y(n3574) );
  NOR2X1 U425 ( .A(n3492), .B(n3493), .Y(n66) );
  NOR2X1 U426 ( .A(n3492), .B(n3503), .Y(n3570) );
  NOR2X1 U427 ( .A(n3496), .B(n3502), .Y(n3566) );
  NOR2X1 U428 ( .A(n3495), .B(n3502), .Y(n3576) );
  NOR2X1 U429 ( .A(n3497), .B(n3502), .Y(n3545) );
  NOR2X1 U430 ( .A(n3496), .B(n3506), .Y(n3564) );
  NOR2X1 U431 ( .A(n3496), .B(n3498), .Y(n3519) );
  NOR2X1 U432 ( .A(n3495), .B(n3506), .Y(n3520) );
  NOR2X1 U433 ( .A(n3495), .B(n3498), .Y(n3542) );
  NOR2X1 U434 ( .A(n3497), .B(n3506), .Y(n3557) );
  NOR2X1 U435 ( .A(n3497), .B(n3498), .Y(n3581) );
  NOR2X1 U436 ( .A(n3496), .B(n3504), .Y(n3540) );
  NOR2X1 U437 ( .A(n3495), .B(n3504), .Y(n3521) );
  NOR2X1 U438 ( .A(n3497), .B(n3504), .Y(n3556) );
  NOR2X1 U439 ( .A(n3496), .B(n3501), .Y(n3522) );
  NOR2X1 U440 ( .A(n3495), .B(n3501), .Y(n3523) );
  NOR2X1 U441 ( .A(n3497), .B(n3501), .Y(n3544) );
  NOR2X1 U442 ( .A(n3496), .B(n3503), .Y(n3541) );
  NOR2X1 U443 ( .A(n3495), .B(n3503), .Y(n3572) );
  NOR2X1 U444 ( .A(n3497), .B(n3503), .Y(n3543) );
  NOR2X1 U445 ( .A(n3499), .B(n3502), .Y(n3561) );
  NOR2X1 U446 ( .A(n3500), .B(n3502), .Y(n3524) );
  NOR2X1 U447 ( .A(n3499), .B(n3506), .Y(n3567) );
  NOR2X1 U448 ( .A(n3500), .B(n3506), .Y(n3531) );
  NOR2X1 U449 ( .A(n3499), .B(n3504), .Y(n3573) );
  NOR2X1 U450 ( .A(n3500), .B(n3504), .Y(n3535) );
  NOR2X1 U451 ( .A(n3499), .B(n3501), .Y(n3577) );
  NOR2X1 U452 ( .A(n3500), .B(n3501), .Y(n3529) );
  NOR2X1 U453 ( .A(n3499), .B(n3503), .Y(n3575) );
  NOR2X1 U454 ( .A(n3500), .B(n3503), .Y(n3539) );
  NOR2X1 U455 ( .A(n3505), .B(n3506), .Y(n3532) );
  CLKINVX3 U456 ( .A(n16075), .Y(n18130) );
  AND2X2 U457 ( .A(n3485), .B(n3491), .Y(n2085) );
  CLKINVX3 U458 ( .A(n16074), .Y(n18129) );
  CLKINVX3 U459 ( .A(n16077), .Y(n18245) );
  CLKINVX3 U460 ( .A(n16076), .Y(n18127) );
  CLKINVX3 U461 ( .A(n18173), .Y(n18167) );
  CLKINVX3 U462 ( .A(n18159), .Y(n18153) );
  INVX1 U463 ( .A(n2083), .Y(n18159) );
  CLKINVX3 U464 ( .A(n18215), .Y(n18209) );
  INVX1 U465 ( .A(n2080), .Y(n18180) );
  INVX1 U466 ( .A(n2086), .Y(n18138) );
  INVX1 U467 ( .A(n2072), .Y(n18208) );
  CLKINVX3 U468 ( .A(n18194), .Y(n18188) );
  INVX1 U469 ( .A(n2079), .Y(n18187) );
  INVX1 U470 ( .A(n2082), .Y(n18166) );
  INVX1 U471 ( .A(n2081), .Y(n18173) );
  INVX1 U472 ( .A(n2084), .Y(n18152) );
  INVX1 U473 ( .A(n2068), .Y(n18236) );
  INVX1 U474 ( .A(n2070), .Y(n18222) );
  INVX1 U475 ( .A(n2069), .Y(n18229) );
  INVX1 U476 ( .A(n2074), .Y(n18194) );
  INVX1 U477 ( .A(n2073), .Y(n18201) );
  INVX1 U478 ( .A(n2067), .Y(n18243) );
  INVX1 U479 ( .A(n2071), .Y(n18215) );
  INVX1 U480 ( .A(\wd<0> ), .Y(n18441) );
  INVX1 U481 ( .A(\wd<1> ), .Y(n18445) );
  INVX1 U482 ( .A(\wd<2> ), .Y(n18449) );
  INVX1 U483 ( .A(\wd<3> ), .Y(n18453) );
  INVX1 U484 ( .A(\wd<4> ), .Y(n18457) );
  INVX1 U485 ( .A(\wd<5> ), .Y(n18461) );
  INVX1 U486 ( .A(\wd<6> ), .Y(n18465) );
  INVX1 U487 ( .A(\wd<7> ), .Y(n18469) );
  INVX1 U488 ( .A(\wd<8> ), .Y(n18473) );
  INVX1 U489 ( .A(\wd<9> ), .Y(n18477) );
  INVX1 U490 ( .A(\wd<10> ), .Y(n18481) );
  INVX1 U491 ( .A(\wd<11> ), .Y(n18485) );
  INVX1 U492 ( .A(\wd<12> ), .Y(n18489) );
  INVX1 U493 ( .A(\wd<13> ), .Y(n18493) );
  INVX1 U494 ( .A(\wd<14> ), .Y(n18497) );
  INVX1 U495 ( .A(\wd<15> ), .Y(n18501) );
  INVX1 U496 ( .A(\wd<16> ), .Y(n18505) );
  INVX1 U497 ( .A(\wd<17> ), .Y(n18509) );
  INVX1 U498 ( .A(\wd<18> ), .Y(n18513) );
  INVX1 U499 ( .A(\wd<19> ), .Y(n18517) );
  INVX1 U500 ( .A(\wd<20> ), .Y(n18521) );
  INVX1 U501 ( .A(\wd<21> ), .Y(n18525) );
  INVX1 U502 ( .A(\wd<22> ), .Y(n18529) );
  INVX1 U503 ( .A(\wd<23> ), .Y(n18533) );
  INVX1 U504 ( .A(\wd<24> ), .Y(n18537) );
  INVX1 U505 ( .A(\wd<25> ), .Y(n18541) );
  INVX1 U506 ( .A(\wd<26> ), .Y(n18545) );
  INVX1 U507 ( .A(\wd<27> ), .Y(n18549) );
  INVX1 U508 ( .A(\wd<28> ), .Y(n18553) );
  INVX1 U509 ( .A(\wd<29> ), .Y(n18557) );
  INVX1 U510 ( .A(\wd<30> ), .Y(n18561) );
  INVX1 U511 ( .A(\wd<31> ), .Y(n18565) );
  NAND2X2 U512 ( .A(n3507), .B(n18126), .Y(n3495) );
  NAND2X2 U513 ( .A(n3507), .B(n18130), .Y(n3497) );
  NAND2X2 U514 ( .A(n3507), .B(n18244), .Y(n3499) );
  NAND2X2 U515 ( .A(n3507), .B(n18128), .Y(n3500) );
  AND2X2 U516 ( .A(n3512), .B(n18568), .Y(n3509) );
  CLKINVX3 U517 ( .A(n16074), .Y(n18128) );
  CLKINVX3 U518 ( .A(n16077), .Y(n18244) );
  CLKINVX3 U519 ( .A(n16076), .Y(n18126) );
  NAND2X2 U520 ( .A(n3510), .B(n3482), .Y(n3494) );
  NAND2X2 U521 ( .A(n3511), .B(n3485), .Y(n3493) );
  NAND2X2 U522 ( .A(n3511), .B(n3481), .Y(n3498) );
  NAND2X2 U523 ( .A(n3511), .B(n3482), .Y(n3502) );
  NAND2X2 U524 ( .A(n3510), .B(n3483), .Y(n3504) );
  NAND2X2 U525 ( .A(n3510), .B(n3485), .Y(n3501) );
  NAND2X2 U526 ( .A(n3511), .B(n3483), .Y(n3503) );
  NAND2X2 U527 ( .A(n3510), .B(n3481), .Y(n3506) );
  NOR2X2 U528 ( .A(n18571), .B(n18570), .Y(n3485) );
  AND2X2 U529 ( .A(n3481), .B(n3490), .Y(n2080) );
  AND2X2 U530 ( .A(n3482), .B(n3490), .Y(n2079) );
  AND2X2 U531 ( .A(n3483), .B(n3490), .Y(n2082) );
  AND2X2 U532 ( .A(n3483), .B(n3491), .Y(n2081) );
  AND2X2 U533 ( .A(n3485), .B(n3490), .Y(n2083) );
  AND2X2 U534 ( .A(n3491), .B(n3482), .Y(n2084) );
  AND2X2 U535 ( .A(n3491), .B(n3481), .Y(n2086) );
  AND2X2 U536 ( .A(n3480), .B(n3481), .Y(n2068) );
  AND2X2 U537 ( .A(n3480), .B(n3482), .Y(n2067) );
  AND2X2 U538 ( .A(n3484), .B(n3482), .Y(n2072) );
  AND2X2 U539 ( .A(n3480), .B(n3485), .Y(n2071) );
  AND2X2 U540 ( .A(n3480), .B(n3483), .Y(n2070) );
  AND2X2 U541 ( .A(n3484), .B(n3483), .Y(n2069) );
  AND2X2 U542 ( .A(n3484), .B(n3481), .Y(n2074) );
  AND2X2 U543 ( .A(n3484), .B(n3485), .Y(n2073) );
  NOR2X1 U544 ( .A(n18569), .B(n18568), .Y(n3491) );
  AND2X2 U545 ( .A(n3512), .B(N35), .Y(n3507) );
  NOR4BX1 U546 ( .AN(n3517), .B(\a<30> ), .C(\a<28> ), .D(\a<29> ), .Y(n3516)
         );
  NOR3X1 U547 ( .A(\a<31> ), .B(\a<9> ), .C(\a<8> ), .Y(n3517) );
  AND4X2 U548 ( .A(n3513), .B(n3514), .C(n3515), .D(n3516), .Y(n3512) );
  NOR4BX1 U549 ( .AN(n3547), .B(\a<12> ), .C(\a<10> ), .D(\a<11> ), .Y(n3513)
         );
  NOR4BX1 U550 ( .AN(n3537), .B(\a<18> ), .C(\a<16> ), .D(\a<17> ), .Y(n3514)
         );
  NOR4BX1 U551 ( .AN(n3518), .B(\a<24> ), .C(\a<22> ), .D(\a<23> ), .Y(n3515)
         );
  NOR3X1 U552 ( .A(\a<25> ), .B(\a<27> ), .C(\a<26> ), .Y(n3518) );
  NOR3X1 U553 ( .A(\a<19> ), .B(\a<21> ), .C(\a<20> ), .Y(n3537) );
  NOR3X1 U554 ( .A(\a<13> ), .B(\a<15> ), .C(\a<14> ), .Y(n3547) );
  INVX1 U555 ( .A(N37), .Y(n18566) );
  NOR2X2 U556 ( .A(N32), .B(N33), .Y(n3481) );
  NOR2X2 U557 ( .A(n18570), .B(N32), .Y(n3482) );
  NOR2X2 U558 ( .A(n18571), .B(N33), .Y(n3483) );
  NOR2X1 U559 ( .A(n18568), .B(N34), .Y(n3490) );
  NOR2X1 U560 ( .A(N34), .B(N35), .Y(n3480) );
  NOR2X1 U561 ( .A(n18569), .B(N35), .Y(n3484) );
  AND2X2 U562 ( .A(we), .B(n18569), .Y(n3510) );
  AND2X2 U563 ( .A(we), .B(N34), .Y(n3511) );
  NAND4X1 U564 ( .A(n2692), .B(n2693), .C(n2694), .D(n2695), .Y(\rd<25> ) );
  OAI21XL U565 ( .A0(n2726), .A1(n2727), .B0(n18127), .Y(n2692) );
  OAI21XL U566 ( .A0(n2706), .A1(n2707), .B0(n18131), .Y(n2694) );
  OAI21XL U567 ( .A0(n2696), .A1(n2697), .B0(n18245), .Y(n2695) );
  NAND4X1 U568 ( .A(n2472), .B(n2473), .C(n2474), .D(n2475), .Y(\rd<2> ) );
  OAI21XL U569 ( .A0(n2506), .A1(n2507), .B0(n18127), .Y(n2472) );
  OAI21XL U570 ( .A0(n2486), .A1(n2487), .B0(n18131), .Y(n2474) );
  OAI21XL U571 ( .A0(n2476), .A1(n2477), .B0(n18245), .Y(n2475) );
  NAND4X1 U572 ( .A(n2340), .B(n2341), .C(n2342), .D(n2343), .Y(\rd<3> ) );
  OAI21XL U573 ( .A0(n2374), .A1(n2375), .B0(n18127), .Y(n2340) );
  OAI21XL U574 ( .A0(n2354), .A1(n2355), .B0(n18131), .Y(n2342) );
  OAI21XL U575 ( .A0(n2344), .A1(n2345), .B0(n18245), .Y(n2343) );
  NAND4X1 U576 ( .A(n2296), .B(n2297), .C(n2298), .D(n2299), .Y(\rd<4> ) );
  OAI21XL U577 ( .A0(n2330), .A1(n2331), .B0(n18127), .Y(n2296) );
  OAI21XL U578 ( .A0(n2310), .A1(n2311), .B0(n18131), .Y(n2298) );
  OAI21XL U579 ( .A0(n2300), .A1(n2301), .B0(n18245), .Y(n2299) );
  NAND4X1 U580 ( .A(n2252), .B(n2253), .C(n2254), .D(n2255), .Y(\rd<5> ) );
  OAI21XL U581 ( .A0(n2286), .A1(n2287), .B0(n18127), .Y(n2252) );
  OAI21XL U582 ( .A0(n2266), .A1(n2267), .B0(n18131), .Y(n2254) );
  OAI21XL U583 ( .A0(n2256), .A1(n2257), .B0(n18245), .Y(n2255) );
  NAND4X1 U584 ( .A(n2208), .B(n2209), .C(n2210), .D(n2211), .Y(\rd<6> ) );
  OAI21XL U585 ( .A0(n2242), .A1(n2243), .B0(n18127), .Y(n2208) );
  OAI21XL U586 ( .A0(n2222), .A1(n2223), .B0(n18131), .Y(n2210) );
  OAI21XL U587 ( .A0(n2212), .A1(n2213), .B0(n18245), .Y(n2211) );
  NAND4X1 U588 ( .A(n2164), .B(n2165), .C(n2166), .D(n2167), .Y(\rd<7> ) );
  OAI21XL U589 ( .A0(n2198), .A1(n2199), .B0(n18127), .Y(n2164) );
  OAI21XL U590 ( .A0(n2178), .A1(n2179), .B0(n18131), .Y(n2166) );
  OAI21XL U591 ( .A0(n2168), .A1(n2169), .B0(n18245), .Y(n2167) );
  NAND4X1 U592 ( .A(n3396), .B(n3397), .C(n3398), .D(n3399), .Y(\rd<10> ) );
  OAI21XL U593 ( .A0(n3430), .A1(n3431), .B0(n18126), .Y(n3396) );
  OAI21XL U594 ( .A0(n3410), .A1(n3411), .B0(n18130), .Y(n3398) );
  OAI21XL U595 ( .A0(n3400), .A1(n3401), .B0(n18244), .Y(n3399) );
  NAND4X1 U596 ( .A(n3352), .B(n3353), .C(n3354), .D(n3355), .Y(\rd<11> ) );
  OAI21XL U597 ( .A0(n3386), .A1(n3387), .B0(n18126), .Y(n3352) );
  OAI21XL U598 ( .A0(n3366), .A1(n3367), .B0(n18130), .Y(n3354) );
  OAI21XL U599 ( .A0(n3356), .A1(n3357), .B0(n18244), .Y(n3355) );
  NAND4X1 U600 ( .A(n3308), .B(n3309), .C(n3310), .D(n3311), .Y(\rd<12> ) );
  OAI21XL U601 ( .A0(n3342), .A1(n3343), .B0(n18126), .Y(n3308) );
  OAI21XL U602 ( .A0(n3322), .A1(n3323), .B0(n18130), .Y(n3310) );
  OAI21XL U603 ( .A0(n3332), .A1(n3333), .B0(n18128), .Y(n3309) );
  NAND4X1 U604 ( .A(n3264), .B(n3265), .C(n3266), .D(n3267), .Y(\rd<13> ) );
  OAI21XL U605 ( .A0(n3298), .A1(n3299), .B0(n18126), .Y(n3264) );
  OAI21XL U606 ( .A0(n3278), .A1(n3279), .B0(n18130), .Y(n3266) );
  OAI21XL U607 ( .A0(n3288), .A1(n3289), .B0(n18128), .Y(n3265) );
  NAND4X1 U608 ( .A(n3220), .B(n3221), .C(n3222), .D(n3223), .Y(\rd<14> ) );
  OAI21XL U609 ( .A0(n3254), .A1(n3255), .B0(n18126), .Y(n3220) );
  OAI21XL U610 ( .A0(n3234), .A1(n3235), .B0(n18130), .Y(n3222) );
  OAI21XL U611 ( .A0(n3244), .A1(n3245), .B0(n18128), .Y(n3221) );
  NAND4X1 U612 ( .A(n3176), .B(n3177), .C(n3178), .D(n3179), .Y(\rd<15> ) );
  OAI21XL U613 ( .A0(n3210), .A1(n3211), .B0(n18126), .Y(n3176) );
  OAI21XL U614 ( .A0(n3190), .A1(n3191), .B0(n18130), .Y(n3178) );
  OAI21XL U615 ( .A0(n3200), .A1(n3201), .B0(n18128), .Y(n3177) );
  NAND4X1 U616 ( .A(n3132), .B(n3133), .C(n3134), .D(n3135), .Y(\rd<16> ) );
  OAI21XL U617 ( .A0(n3166), .A1(n3167), .B0(n18126), .Y(n3132) );
  OAI21XL U618 ( .A0(n3146), .A1(n3147), .B0(n18130), .Y(n3134) );
  OAI21XL U619 ( .A0(n3136), .A1(n3137), .B0(n18244), .Y(n3135) );
  NAND4X1 U620 ( .A(n3088), .B(n3089), .C(n3090), .D(n3091), .Y(\rd<17> ) );
  OAI21XL U621 ( .A0(n3122), .A1(n3123), .B0(n18126), .Y(n3088) );
  OAI21XL U622 ( .A0(n3102), .A1(n3103), .B0(n18130), .Y(n3090) );
  OAI21XL U623 ( .A0(n3092), .A1(n3093), .B0(n18244), .Y(n3091) );
  NAND4X1 U624 ( .A(n3044), .B(n3045), .C(n3046), .D(n3047), .Y(\rd<18> ) );
  OAI21XL U625 ( .A0(n3078), .A1(n3079), .B0(n18126), .Y(n3044) );
  OAI21XL U626 ( .A0(n3058), .A1(n3059), .B0(n18130), .Y(n3046) );
  OAI21XL U627 ( .A0(n3048), .A1(n3049), .B0(n18244), .Y(n3047) );
  NAND4X1 U628 ( .A(n3000), .B(n3001), .C(n3002), .D(n3003), .Y(\rd<19> ) );
  OAI21XL U629 ( .A0(n3034), .A1(n3035), .B0(n18126), .Y(n3000) );
  OAI21XL U630 ( .A0(n3014), .A1(n3015), .B0(n18130), .Y(n3002) );
  OAI21XL U631 ( .A0(n3004), .A1(n3005), .B0(n18244), .Y(n3003) );
  NAND4X1 U632 ( .A(n2120), .B(n2121), .C(n2122), .D(n2123), .Y(\rd<8> ) );
  OAI21XL U633 ( .A0(n2154), .A1(n2155), .B0(n18127), .Y(n2120) );
  OAI21XL U634 ( .A0(n2134), .A1(n2135), .B0(n18131), .Y(n2122) );
  OAI21XL U635 ( .A0(n2124), .A1(n2125), .B0(n18245), .Y(n2123) );
  NAND4X1 U636 ( .A(n2056), .B(n2057), .C(n2058), .D(n2059), .Y(\rd<9> ) );
  OAI21XL U637 ( .A0(n2109), .A1(n2110), .B0(n18127), .Y(n2056) );
  OAI21XL U638 ( .A0(n2087), .A1(n2088), .B0(n18131), .Y(n2058) );
  OAI21XL U639 ( .A0(n2060), .A1(n2061), .B0(n18245), .Y(n2059) );
  NAND4X1 U640 ( .A(n2912), .B(n2913), .C(n2914), .D(n2915), .Y(\rd<20> ) );
  OAI21XL U641 ( .A0(n2946), .A1(n2947), .B0(n18127), .Y(n2912) );
  OAI21XL U642 ( .A0(n2926), .A1(n2927), .B0(n18131), .Y(n2914) );
  OAI21XL U643 ( .A0(n2936), .A1(n2937), .B0(n18129), .Y(n2913) );
  NAND4X1 U644 ( .A(n2868), .B(n2869), .C(n2870), .D(n2871), .Y(\rd<21> ) );
  OAI21XL U645 ( .A0(n2902), .A1(n2903), .B0(n18127), .Y(n2868) );
  OAI21XL U646 ( .A0(n2882), .A1(n2883), .B0(n18131), .Y(n2870) );
  OAI21XL U647 ( .A0(n2872), .A1(n2873), .B0(n18245), .Y(n2871) );
  NAND4X1 U648 ( .A(n2824), .B(n2825), .C(n2826), .D(n2827), .Y(\rd<22> ) );
  OAI21XL U649 ( .A0(n2858), .A1(n2859), .B0(n18127), .Y(n2824) );
  OAI21XL U650 ( .A0(n2838), .A1(n2839), .B0(n18131), .Y(n2826) );
  OAI21XL U651 ( .A0(n2828), .A1(n2829), .B0(n18245), .Y(n2827) );
  NAND4X1 U652 ( .A(n2780), .B(n2781), .C(n2782), .D(n2783), .Y(\rd<23> ) );
  OAI21XL U653 ( .A0(n2814), .A1(n2815), .B0(n18127), .Y(n2780) );
  OAI21XL U654 ( .A0(n2794), .A1(n2795), .B0(n18131), .Y(n2782) );
  OAI21XL U655 ( .A0(n2784), .A1(n2785), .B0(n18245), .Y(n2783) );
  NAND4X1 U656 ( .A(n2736), .B(n2737), .C(n2738), .D(n2739), .Y(\rd<24> ) );
  OAI21XL U657 ( .A0(n2770), .A1(n2771), .B0(n18127), .Y(n2736) );
  OAI21XL U658 ( .A0(n2750), .A1(n2751), .B0(n18131), .Y(n2738) );
  OAI21XL U659 ( .A0(n2740), .A1(n2741), .B0(n18245), .Y(n2739) );
  NAND4X1 U660 ( .A(n2648), .B(n2649), .C(n2650), .D(n2651), .Y(\rd<26> ) );
  OAI21XL U661 ( .A0(n2682), .A1(n2683), .B0(n18127), .Y(n2648) );
  OAI21XL U662 ( .A0(n2662), .A1(n2663), .B0(n18131), .Y(n2650) );
  OAI21XL U663 ( .A0(n2672), .A1(n2673), .B0(n18129), .Y(n2649) );
  NAND4X1 U664 ( .A(n2604), .B(n2605), .C(n2606), .D(n2607), .Y(\rd<27> ) );
  OAI21XL U665 ( .A0(n2638), .A1(n2639), .B0(n18127), .Y(n2604) );
  OAI21XL U666 ( .A0(n2618), .A1(n2619), .B0(n18131), .Y(n2606) );
  OAI21XL U667 ( .A0(n2628), .A1(n2629), .B0(n18129), .Y(n2605) );
  NAND4X1 U668 ( .A(n2560), .B(n2561), .C(n2562), .D(n2563), .Y(\rd<28> ) );
  OAI21XL U669 ( .A0(n2594), .A1(n2595), .B0(n18127), .Y(n2560) );
  OAI21XL U670 ( .A0(n2584), .A1(n2585), .B0(n18129), .Y(n2561) );
  OAI21XL U671 ( .A0(n2574), .A1(n2575), .B0(n18131), .Y(n2562) );
  NAND4X1 U672 ( .A(n2516), .B(n2517), .C(n2518), .D(n2519), .Y(\rd<29> ) );
  OAI21XL U673 ( .A0(n2550), .A1(n2551), .B0(n18127), .Y(n2516) );
  OAI21XL U674 ( .A0(n2540), .A1(n2541), .B0(n18129), .Y(n2517) );
  OAI21XL U675 ( .A0(n2530), .A1(n2531), .B0(n18131), .Y(n2518) );
  NAND4X1 U676 ( .A(n2428), .B(n2429), .C(n2430), .D(n2431), .Y(\rd<30> ) );
  OAI21XL U677 ( .A0(n2462), .A1(n2463), .B0(n18127), .Y(n2428) );
  OAI21XL U678 ( .A0(n2442), .A1(n2443), .B0(n18131), .Y(n2430) );
  OAI21XL U679 ( .A0(n2452), .A1(n2453), .B0(n18129), .Y(n2429) );
  NAND4X1 U680 ( .A(n2384), .B(n2385), .C(n2386), .D(n2387), .Y(\rd<31> ) );
  OAI21XL U681 ( .A0(n2418), .A1(n2419), .B0(n18127), .Y(n2384) );
  OAI21XL U682 ( .A0(n2398), .A1(n2399), .B0(n18131), .Y(n2386) );
  OAI21XL U683 ( .A0(n2388), .A1(n2389), .B0(n18245), .Y(n2387) );
  NAND4X1 U684 ( .A(n3440), .B(n3441), .C(n3442), .D(n3443), .Y(\rd<0> ) );
  OAI21XL U685 ( .A0(n3474), .A1(n3475), .B0(n18126), .Y(n3440) );
  OAI21XL U686 ( .A0(n3454), .A1(n3455), .B0(n18130), .Y(n3442) );
  OAI21XL U687 ( .A0(n3444), .A1(n3445), .B0(n18244), .Y(n3443) );
  NAND4X1 U688 ( .A(n2956), .B(n2957), .C(n2958), .D(n2959), .Y(\rd<1> ) );
  OAI21XL U689 ( .A0(n2990), .A1(n2991), .B0(n18127), .Y(n2956) );
  OAI21XL U690 ( .A0(n2970), .A1(n2971), .B0(n18131), .Y(n2958) );
  OAI21XL U691 ( .A0(n2960), .A1(n2961), .B0(n18245), .Y(n2959) );
  INVX1 U692 ( .A(N34), .Y(n18569) );
  INVX1 U693 ( .A(N35), .Y(n18568) );
  INVX1 U694 ( .A(N32), .Y(n18571) );
  INVX1 U695 ( .A(N36), .Y(n18567) );
  INVX1 U696 ( .A(N33), .Y(n18570) );
  AOI22X1 U697 ( .A0(n18186), .A1(\RAM<42><2> ), .B0(n18175), .B1(\RAM<40><2> ), .Y(n2505) );
  AOI22X1 U698 ( .A0(n18241), .A1(\RAM<34><2> ), .B0(n18234), .B1(\RAM<32><2> ), .Y(n2501) );
  AOI22X1 U699 ( .A0(n18183), .A1(\RAM<10><2> ), .B0(n18177), .B1(\RAM<8><2> ), 
        .Y(n2485) );
  AOI22X1 U700 ( .A0(n2067), .A1(\RAM<2><2> ), .B0(n18234), .B1(\RAM<0><2> ), 
        .Y(n2481) );
  AOI22X1 U701 ( .A0(n18186), .A1(\RAM<58><2> ), .B0(n18175), .B1(\RAM<56><2> ), .Y(n2495) );
  AOI22X1 U702 ( .A0(n18239), .A1(\RAM<50><2> ), .B0(n18234), .B1(\RAM<48><2> ), .Y(n2491) );
  AOI22X1 U703 ( .A0(n18181), .A1(\RAM<26><2> ), .B0(n18175), .B1(\RAM<24><2> ), .Y(n2515) );
  AOI22X1 U704 ( .A0(n18240), .A1(\RAM<18><2> ), .B0(n18234), .B1(\RAM<16><2> ), .Y(n2511) );
  AOI22X1 U705 ( .A0(n18185), .A1(\RAM<42><3> ), .B0(n18178), .B1(\RAM<40><3> ), .Y(n2373) );
  AOI22X1 U706 ( .A0(n18241), .A1(\RAM<34><3> ), .B0(n18232), .B1(\RAM<32><3> ), .Y(n2369) );
  AOI22X1 U707 ( .A0(n18185), .A1(\RAM<10><3> ), .B0(n18178), .B1(\RAM<8><3> ), 
        .Y(n2353) );
  AOI22X1 U708 ( .A0(n18241), .A1(\RAM<2><3> ), .B0(n18232), .B1(\RAM<0><3> ), 
        .Y(n2349) );
  AOI22X1 U709 ( .A0(n18185), .A1(\RAM<58><3> ), .B0(n18178), .B1(\RAM<56><3> ), .Y(n2363) );
  AOI22X1 U710 ( .A0(n18241), .A1(\RAM<50><3> ), .B0(n18232), .B1(\RAM<48><3> ), .Y(n2359) );
  AOI22X1 U711 ( .A0(n18185), .A1(\RAM<26><3> ), .B0(n18178), .B1(\RAM<24><3> ), .Y(n2383) );
  AOI22X1 U712 ( .A0(n18241), .A1(\RAM<18><3> ), .B0(n18232), .B1(\RAM<16><3> ), .Y(n2379) );
  AOI22X1 U713 ( .A0(n18185), .A1(\RAM<42><4> ), .B0(n18178), .B1(\RAM<40><4> ), .Y(n2329) );
  AOI22X1 U714 ( .A0(n18241), .A1(\RAM<34><4> ), .B0(n18234), .B1(\RAM<32><4> ), .Y(n2325) );
  AOI22X1 U715 ( .A0(n18185), .A1(\RAM<10><4> ), .B0(n18178), .B1(\RAM<8><4> ), 
        .Y(n2309) );
  AOI22X1 U716 ( .A0(n18241), .A1(\RAM<2><4> ), .B0(n18234), .B1(\RAM<0><4> ), 
        .Y(n2305) );
  AOI22X1 U717 ( .A0(n18185), .A1(\RAM<58><4> ), .B0(n18178), .B1(\RAM<56><4> ), .Y(n2319) );
  AOI22X1 U718 ( .A0(n18241), .A1(\RAM<50><4> ), .B0(n18234), .B1(\RAM<48><4> ), .Y(n2315) );
  AOI22X1 U719 ( .A0(n18185), .A1(\RAM<26><4> ), .B0(n18178), .B1(\RAM<24><4> ), .Y(n2339) );
  AOI22X1 U720 ( .A0(n18241), .A1(\RAM<18><4> ), .B0(n18234), .B1(\RAM<16><4> ), .Y(n2335) );
  AOI22X1 U721 ( .A0(n18186), .A1(\RAM<42><5> ), .B0(n18179), .B1(\RAM<40><5> ), .Y(n2285) );
  AOI22X1 U722 ( .A0(n18242), .A1(\RAM<34><5> ), .B0(n18235), .B1(\RAM<32><5> ), .Y(n2281) );
  AOI22X1 U723 ( .A0(n18186), .A1(\RAM<10><5> ), .B0(n18179), .B1(\RAM<8><5> ), 
        .Y(n2265) );
  AOI22X1 U724 ( .A0(n18242), .A1(\RAM<2><5> ), .B0(n18235), .B1(\RAM<0><5> ), 
        .Y(n2261) );
  AOI22X1 U725 ( .A0(n18186), .A1(\RAM<58><5> ), .B0(n18179), .B1(\RAM<56><5> ), .Y(n2275) );
  AOI22X1 U726 ( .A0(n18242), .A1(\RAM<50><5> ), .B0(n18235), .B1(\RAM<48><5> ), .Y(n2271) );
  AOI22X1 U727 ( .A0(n18186), .A1(\RAM<26><5> ), .B0(n18179), .B1(\RAM<24><5> ), .Y(n2295) );
  AOI22X1 U728 ( .A0(n18242), .A1(\RAM<18><5> ), .B0(n18235), .B1(\RAM<16><5> ), .Y(n2291) );
  AOI22X1 U729 ( .A0(n18186), .A1(\RAM<42><6> ), .B0(n18179), .B1(\RAM<40><6> ), .Y(n2241) );
  AOI22X1 U730 ( .A0(n18242), .A1(\RAM<34><6> ), .B0(n18235), .B1(\RAM<32><6> ), .Y(n2237) );
  AOI22X1 U731 ( .A0(n18186), .A1(\RAM<10><6> ), .B0(n18179), .B1(\RAM<8><6> ), 
        .Y(n2221) );
  AOI22X1 U732 ( .A0(n18242), .A1(\RAM<2><6> ), .B0(n18235), .B1(\RAM<0><6> ), 
        .Y(n2217) );
  AOI22X1 U733 ( .A0(n18186), .A1(\RAM<58><6> ), .B0(n18179), .B1(\RAM<56><6> ), .Y(n2231) );
  AOI22X1 U734 ( .A0(n18242), .A1(\RAM<50><6> ), .B0(n18235), .B1(\RAM<48><6> ), .Y(n2227) );
  AOI22X1 U735 ( .A0(n18186), .A1(\RAM<26><6> ), .B0(n18179), .B1(\RAM<24><6> ), .Y(n2251) );
  AOI22X1 U736 ( .A0(n18242), .A1(\RAM<18><6> ), .B0(n18235), .B1(\RAM<16><6> ), .Y(n2247) );
  AOI22X1 U737 ( .A0(n18186), .A1(\RAM<42><7> ), .B0(n18179), .B1(\RAM<40><7> ), .Y(n2197) );
  AOI22X1 U738 ( .A0(n18242), .A1(\RAM<34><7> ), .B0(n18235), .B1(\RAM<32><7> ), .Y(n2193) );
  AOI22X1 U739 ( .A0(n18186), .A1(\RAM<10><7> ), .B0(n18179), .B1(\RAM<8><7> ), 
        .Y(n2177) );
  AOI22X1 U740 ( .A0(n18242), .A1(\RAM<2><7> ), .B0(n18235), .B1(\RAM<0><7> ), 
        .Y(n2173) );
  AOI22X1 U741 ( .A0(n18186), .A1(\RAM<58><7> ), .B0(n18179), .B1(\RAM<56><7> ), .Y(n2187) );
  AOI22X1 U742 ( .A0(n18242), .A1(\RAM<50><7> ), .B0(n18235), .B1(\RAM<48><7> ), .Y(n2183) );
  AOI22X1 U743 ( .A0(n18186), .A1(\RAM<26><7> ), .B0(n18179), .B1(\RAM<24><7> ), .Y(n2207) );
  AOI22X1 U744 ( .A0(n18242), .A1(\RAM<18><7> ), .B0(n18235), .B1(\RAM<16><7> ), .Y(n2203) );
  AOI22X1 U745 ( .A0(n18185), .A1(\RAM<42><8> ), .B0(n18178), .B1(\RAM<40><8> ), .Y(n2153) );
  AOI22X1 U746 ( .A0(n18237), .A1(\RAM<34><8> ), .B0(n18234), .B1(\RAM<32><8> ), .Y(n2149) );
  AOI22X1 U747 ( .A0(n2079), .A1(\RAM<10><8> ), .B0(n18179), .B1(\RAM<8><8> ), 
        .Y(n2133) );
  AOI22X1 U748 ( .A0(n18241), .A1(\RAM<2><8> ), .B0(n18232), .B1(\RAM<0><8> ), 
        .Y(n2129) );
  AOI22X1 U749 ( .A0(n18184), .A1(\RAM<58><8> ), .B0(n18177), .B1(\RAM<56><8> ), .Y(n2143) );
  AOI22X1 U750 ( .A0(n18238), .A1(\RAM<50><8> ), .B0(n18233), .B1(\RAM<48><8> ), .Y(n2139) );
  AOI22X1 U751 ( .A0(n18183), .A1(\RAM<26><8> ), .B0(n18179), .B1(\RAM<24><8> ), .Y(n2163) );
  AOI22X1 U752 ( .A0(n18238), .A1(\RAM<18><8> ), .B0(n18232), .B1(\RAM<16><8> ), .Y(n2159) );
  AOI22X1 U753 ( .A0(n18182), .A1(\RAM<42><9> ), .B0(n18178), .B1(\RAM<40><9> ), .Y(n2108) );
  AOI22X1 U754 ( .A0(n18242), .A1(\RAM<34><9> ), .B0(n18235), .B1(\RAM<32><9> ), .Y(n2104) );
  AOI22X1 U755 ( .A0(n2079), .A1(\RAM<10><9> ), .B0(n18176), .B1(\RAM<8><9> ), 
        .Y(n2078) );
  AOI22X1 U756 ( .A0(n2067), .A1(\RAM<2><9> ), .B0(n18235), .B1(\RAM<0><9> ), 
        .Y(n2066) );
  AOI22X1 U757 ( .A0(n2079), .A1(\RAM<58><9> ), .B0(n18176), .B1(\RAM<56><9> ), 
        .Y(n2097) );
  AOI22X1 U758 ( .A0(n18242), .A1(\RAM<50><9> ), .B0(n18235), .B1(\RAM<48><9> ), .Y(n2093) );
  AOI22X1 U759 ( .A0(n18183), .A1(\RAM<26><9> ), .B0(n18179), .B1(\RAM<24><9> ), .Y(n2119) );
  AOI22X1 U760 ( .A0(n18242), .A1(\RAM<18><9> ), .B0(n18235), .B1(\RAM<16><9> ), .Y(n2115) );
  AOI22X1 U761 ( .A0(n18183), .A1(\RAM<42><10> ), .B0(n18178), .B1(
        \RAM<40><10> ), .Y(n3429) );
  AOI22X1 U762 ( .A0(n18238), .A1(\RAM<34><10> ), .B0(n18232), .B1(
        \RAM<32><10> ), .Y(n3425) );
  AOI22X1 U763 ( .A0(n18182), .A1(\RAM<10><10> ), .B0(n18178), .B1(
        \RAM<8><10> ), .Y(n3409) );
  AOI22X1 U764 ( .A0(n18239), .A1(\RAM<2><10> ), .B0(n2068), .B1(\RAM<0><10> ), 
        .Y(n3405) );
  AOI22X1 U765 ( .A0(n18183), .A1(\RAM<58><10> ), .B0(n18179), .B1(
        \RAM<56><10> ), .Y(n3419) );
  AOI22X1 U766 ( .A0(n18238), .A1(\RAM<50><10> ), .B0(n18232), .B1(
        \RAM<48><10> ), .Y(n3415) );
  AOI22X1 U767 ( .A0(n18185), .A1(\RAM<26><10> ), .B0(n18178), .B1(
        \RAM<24><10> ), .Y(n3439) );
  AOI22X1 U768 ( .A0(n18242), .A1(\RAM<18><10> ), .B0(n18232), .B1(
        \RAM<16><10> ), .Y(n3435) );
  AOI22X1 U769 ( .A0(n18185), .A1(\RAM<42><11> ), .B0(n18176), .B1(
        \RAM<40><11> ), .Y(n3385) );
  AOI22X1 U770 ( .A0(n18240), .A1(\RAM<34><11> ), .B0(n18234), .B1(
        \RAM<32><11> ), .Y(n3381) );
  AOI22X1 U771 ( .A0(n2079), .A1(\RAM<10><11> ), .B0(n2080), .B1(\RAM<8><11> ), 
        .Y(n3365) );
  AOI22X1 U772 ( .A0(n2067), .A1(\RAM<2><11> ), .B0(n18233), .B1(\RAM<0><11> ), 
        .Y(n3361) );
  AOI22X1 U773 ( .A0(n18183), .A1(\RAM<58><11> ), .B0(n18178), .B1(
        \RAM<56><11> ), .Y(n3375) );
  AOI22X1 U774 ( .A0(n18241), .A1(\RAM<50><11> ), .B0(n18233), .B1(
        \RAM<48><11> ), .Y(n3371) );
  AOI22X1 U775 ( .A0(n18182), .A1(\RAM<26><11> ), .B0(n18176), .B1(
        \RAM<24><11> ), .Y(n3395) );
  AOI22X1 U776 ( .A0(n18237), .A1(\RAM<18><11> ), .B0(n18234), .B1(
        \RAM<16><11> ), .Y(n3391) );
  AOI22X1 U777 ( .A0(n18181), .A1(\RAM<10><12> ), .B0(n18174), .B1(
        \RAM<8><12> ), .Y(n3321) );
  AOI22X1 U778 ( .A0(n18237), .A1(\RAM<2><12> ), .B0(n18230), .B1(\RAM<0><12> ), .Y(n3317) );
  AOI22X1 U779 ( .A0(n18181), .A1(\RAM<42><12> ), .B0(n18174), .B1(
        \RAM<40><12> ), .Y(n3341) );
  AOI22X1 U780 ( .A0(n18237), .A1(\RAM<34><12> ), .B0(n18230), .B1(
        \RAM<32><12> ), .Y(n3337) );
  AOI22X1 U781 ( .A0(n18181), .A1(\RAM<58><12> ), .B0(n18174), .B1(
        \RAM<56><12> ), .Y(n3331) );
  AOI22X1 U782 ( .A0(n18237), .A1(\RAM<50><12> ), .B0(n18230), .B1(
        \RAM<48><12> ), .Y(n3327) );
  AOI22X1 U783 ( .A0(n18181), .A1(\RAM<26><12> ), .B0(n18174), .B1(
        \RAM<24><12> ), .Y(n3351) );
  AOI22X1 U784 ( .A0(n18237), .A1(\RAM<18><12> ), .B0(n18230), .B1(
        \RAM<16><12> ), .Y(n3347) );
  AOI22X1 U785 ( .A0(n18181), .A1(\RAM<10><13> ), .B0(n18174), .B1(
        \RAM<8><13> ), .Y(n3277) );
  AOI22X1 U786 ( .A0(n18237), .A1(\RAM<2><13> ), .B0(n18230), .B1(\RAM<0><13> ), .Y(n3273) );
  AOI22X1 U787 ( .A0(n18181), .A1(\RAM<42><13> ), .B0(n18174), .B1(
        \RAM<40><13> ), .Y(n3297) );
  AOI22X1 U788 ( .A0(n18237), .A1(\RAM<34><13> ), .B0(n18230), .B1(
        \RAM<32><13> ), .Y(n3293) );
  AOI22X1 U789 ( .A0(n18181), .A1(\RAM<58><13> ), .B0(n18174), .B1(
        \RAM<56><13> ), .Y(n3287) );
  AOI22X1 U790 ( .A0(n18237), .A1(\RAM<50><13> ), .B0(n18230), .B1(
        \RAM<48><13> ), .Y(n3283) );
  AOI22X1 U791 ( .A0(n18181), .A1(\RAM<26><13> ), .B0(n18174), .B1(
        \RAM<24><13> ), .Y(n3307) );
  AOI22X1 U792 ( .A0(n18237), .A1(\RAM<18><13> ), .B0(n18230), .B1(
        \RAM<16><13> ), .Y(n3303) );
  AOI22X1 U793 ( .A0(n18181), .A1(\RAM<10><14> ), .B0(n18174), .B1(
        \RAM<8><14> ), .Y(n3233) );
  AOI22X1 U794 ( .A0(n18237), .A1(\RAM<2><14> ), .B0(n18230), .B1(\RAM<0><14> ), .Y(n3229) );
  AOI22X1 U795 ( .A0(n18181), .A1(\RAM<42><14> ), .B0(n18174), .B1(
        \RAM<40><14> ), .Y(n3253) );
  AOI22X1 U796 ( .A0(n18237), .A1(\RAM<34><14> ), .B0(n18230), .B1(
        \RAM<32><14> ), .Y(n3249) );
  AOI22X1 U797 ( .A0(n18181), .A1(\RAM<58><14> ), .B0(n18174), .B1(
        \RAM<56><14> ), .Y(n3243) );
  AOI22X1 U798 ( .A0(n18237), .A1(\RAM<50><14> ), .B0(n18230), .B1(
        \RAM<48><14> ), .Y(n3239) );
  AOI22X1 U799 ( .A0(n18181), .A1(\RAM<26><14> ), .B0(n18174), .B1(
        \RAM<24><14> ), .Y(n3263) );
  AOI22X1 U800 ( .A0(n18237), .A1(\RAM<18><14> ), .B0(n18230), .B1(
        \RAM<16><14> ), .Y(n3259) );
  AOI22X1 U801 ( .A0(n18182), .A1(\RAM<10><15> ), .B0(n18175), .B1(
        \RAM<8><15> ), .Y(n3189) );
  AOI22X1 U802 ( .A0(n18237), .A1(\RAM<2><15> ), .B0(n18231), .B1(\RAM<0><15> ), .Y(n3185) );
  AOI22X1 U803 ( .A0(n18182), .A1(\RAM<42><15> ), .B0(n18175), .B1(
        \RAM<40><15> ), .Y(n3209) );
  AOI22X1 U804 ( .A0(n18242), .A1(\RAM<34><15> ), .B0(n18231), .B1(
        \RAM<32><15> ), .Y(n3205) );
  AOI22X1 U805 ( .A0(n18182), .A1(\RAM<58><15> ), .B0(n18175), .B1(
        \RAM<56><15> ), .Y(n3199) );
  AOI22X1 U806 ( .A0(n18238), .A1(\RAM<50><15> ), .B0(n18231), .B1(
        \RAM<48><15> ), .Y(n3195) );
  AOI22X1 U807 ( .A0(n18182), .A1(\RAM<26><15> ), .B0(n18175), .B1(
        \RAM<24><15> ), .Y(n3219) );
  AOI22X1 U808 ( .A0(n18237), .A1(\RAM<18><15> ), .B0(n18231), .B1(
        \RAM<16><15> ), .Y(n3215) );
  AOI22X1 U809 ( .A0(n18182), .A1(\RAM<42><16> ), .B0(n18175), .B1(
        \RAM<40><16> ), .Y(n3165) );
  AOI22X1 U810 ( .A0(n18237), .A1(\RAM<34><16> ), .B0(n18231), .B1(
        \RAM<32><16> ), .Y(n3161) );
  AOI22X1 U811 ( .A0(n18182), .A1(\RAM<10><16> ), .B0(n18175), .B1(
        \RAM<8><16> ), .Y(n3145) );
  AOI22X1 U812 ( .A0(n18238), .A1(\RAM<2><16> ), .B0(n18231), .B1(\RAM<0><16> ), .Y(n3141) );
  AOI22X1 U813 ( .A0(n18182), .A1(\RAM<58><16> ), .B0(n18175), .B1(
        \RAM<56><16> ), .Y(n3155) );
  AOI22X1 U814 ( .A0(n18242), .A1(\RAM<50><16> ), .B0(n18231), .B1(
        \RAM<48><16> ), .Y(n3151) );
  AOI22X1 U815 ( .A0(n18182), .A1(\RAM<26><16> ), .B0(n18175), .B1(
        \RAM<24><16> ), .Y(n3175) );
  AOI22X1 U816 ( .A0(n18237), .A1(\RAM<18><16> ), .B0(n18231), .B1(
        \RAM<16><16> ), .Y(n3171) );
  AOI22X1 U817 ( .A0(n18182), .A1(\RAM<42><17> ), .B0(n18175), .B1(
        \RAM<40><17> ), .Y(n3121) );
  AOI22X1 U818 ( .A0(n18237), .A1(\RAM<34><17> ), .B0(n18231), .B1(
        \RAM<32><17> ), .Y(n3117) );
  AOI22X1 U819 ( .A0(n18182), .A1(\RAM<10><17> ), .B0(n18175), .B1(
        \RAM<8><17> ), .Y(n3101) );
  AOI22X1 U820 ( .A0(n18242), .A1(\RAM<2><17> ), .B0(n18231), .B1(\RAM<0><17> ), .Y(n3097) );
  AOI22X1 U821 ( .A0(n18182), .A1(\RAM<58><17> ), .B0(n18175), .B1(
        \RAM<56><17> ), .Y(n3111) );
  AOI22X1 U822 ( .A0(n18237), .A1(\RAM<50><17> ), .B0(n18231), .B1(
        \RAM<48><17> ), .Y(n3107) );
  AOI22X1 U823 ( .A0(n18182), .A1(\RAM<26><17> ), .B0(n18175), .B1(
        \RAM<24><17> ), .Y(n3131) );
  AOI22X1 U824 ( .A0(n18238), .A1(\RAM<18><17> ), .B0(n18231), .B1(
        \RAM<16><17> ), .Y(n3127) );
  AOI22X1 U825 ( .A0(n18184), .A1(\RAM<42><18> ), .B0(n18178), .B1(
        \RAM<40><18> ), .Y(n3077) );
  AOI22X1 U826 ( .A0(n18238), .A1(\RAM<34><18> ), .B0(n18231), .B1(
        \RAM<32><18> ), .Y(n3073) );
  AOI22X1 U827 ( .A0(n18184), .A1(\RAM<10><18> ), .B0(n18174), .B1(
        \RAM<8><18> ), .Y(n3057) );
  AOI22X1 U828 ( .A0(n18238), .A1(\RAM<2><18> ), .B0(n18231), .B1(\RAM<0><18> ), .Y(n3053) );
  AOI22X1 U829 ( .A0(n18181), .A1(\RAM<58><18> ), .B0(n18179), .B1(
        \RAM<56><18> ), .Y(n3067) );
  AOI22X1 U830 ( .A0(n18238), .A1(\RAM<50><18> ), .B0(n18231), .B1(
        \RAM<48><18> ), .Y(n3063) );
  AOI22X1 U831 ( .A0(n18186), .A1(\RAM<26><18> ), .B0(n18178), .B1(
        \RAM<24><18> ), .Y(n3087) );
  AOI22X1 U832 ( .A0(n18238), .A1(\RAM<18><18> ), .B0(n18231), .B1(
        \RAM<16><18> ), .Y(n3083) );
  AOI22X1 U833 ( .A0(n18186), .A1(\RAM<42><19> ), .B0(n18176), .B1(
        \RAM<40><19> ), .Y(n3033) );
  AOI22X1 U834 ( .A0(n18238), .A1(\RAM<34><19> ), .B0(n18230), .B1(
        \RAM<32><19> ), .Y(n3029) );
  AOI22X1 U835 ( .A0(n18181), .A1(\RAM<10><19> ), .B0(n18177), .B1(
        \RAM<8><19> ), .Y(n3013) );
  AOI22X1 U836 ( .A0(n18238), .A1(\RAM<2><19> ), .B0(n18230), .B1(\RAM<0><19> ), .Y(n3009) );
  AOI22X1 U837 ( .A0(n18186), .A1(\RAM<58><19> ), .B0(n18179), .B1(
        \RAM<56><19> ), .Y(n3023) );
  AOI22X1 U838 ( .A0(n18238), .A1(\RAM<50><19> ), .B0(n18230), .B1(
        \RAM<48><19> ), .Y(n3019) );
  AOI22X1 U839 ( .A0(n18186), .A1(\RAM<26><19> ), .B0(n18176), .B1(
        \RAM<24><19> ), .Y(n3043) );
  AOI22X1 U840 ( .A0(n18238), .A1(\RAM<18><19> ), .B0(n18230), .B1(
        \RAM<16><19> ), .Y(n3039) );
  AOI22X1 U841 ( .A0(n18183), .A1(\RAM<10><20> ), .B0(n18176), .B1(
        \RAM<8><20> ), .Y(n2925) );
  AOI22X1 U842 ( .A0(n18239), .A1(\RAM<2><20> ), .B0(n18232), .B1(\RAM<0><20> ), .Y(n2921) );
  AOI22X1 U843 ( .A0(n18183), .A1(\RAM<42><20> ), .B0(n18176), .B1(
        \RAM<40><20> ), .Y(n2945) );
  AOI22X1 U844 ( .A0(n18239), .A1(\RAM<34><20> ), .B0(n18232), .B1(
        \RAM<32><20> ), .Y(n2941) );
  AOI22X1 U845 ( .A0(n18183), .A1(\RAM<58><20> ), .B0(n18176), .B1(
        \RAM<56><20> ), .Y(n2935) );
  AOI22X1 U846 ( .A0(n18239), .A1(\RAM<50><20> ), .B0(n18232), .B1(
        \RAM<48><20> ), .Y(n2931) );
  AOI22X1 U847 ( .A0(n18183), .A1(\RAM<26><20> ), .B0(n18176), .B1(
        \RAM<24><20> ), .Y(n2955) );
  AOI22X1 U848 ( .A0(n18239), .A1(\RAM<18><20> ), .B0(n18232), .B1(
        \RAM<16><20> ), .Y(n2951) );
  AOI22X1 U849 ( .A0(n18183), .A1(\RAM<42><21> ), .B0(n18176), .B1(
        \RAM<40><21> ), .Y(n2901) );
  AOI22X1 U850 ( .A0(n18239), .A1(\RAM<34><21> ), .B0(n18232), .B1(
        \RAM<32><21> ), .Y(n2897) );
  AOI22X1 U851 ( .A0(n18183), .A1(\RAM<10><21> ), .B0(n18176), .B1(
        \RAM<8><21> ), .Y(n2881) );
  AOI22X1 U852 ( .A0(n18239), .A1(\RAM<2><21> ), .B0(n18232), .B1(\RAM<0><21> ), .Y(n2877) );
  AOI22X1 U853 ( .A0(n18183), .A1(\RAM<58><21> ), .B0(n18176), .B1(
        \RAM<56><21> ), .Y(n2891) );
  AOI22X1 U854 ( .A0(n18239), .A1(\RAM<50><21> ), .B0(n18232), .B1(
        \RAM<48><21> ), .Y(n2887) );
  AOI22X1 U855 ( .A0(n18183), .A1(\RAM<26><21> ), .B0(n18176), .B1(
        \RAM<24><21> ), .Y(n2911) );
  AOI22X1 U856 ( .A0(n18239), .A1(\RAM<18><21> ), .B0(n18232), .B1(
        \RAM<16><21> ), .Y(n2907) );
  AOI22X1 U857 ( .A0(n18183), .A1(\RAM<42><22> ), .B0(n18176), .B1(
        \RAM<40><22> ), .Y(n2857) );
  AOI22X1 U858 ( .A0(n18239), .A1(\RAM<34><22> ), .B0(n18232), .B1(
        \RAM<32><22> ), .Y(n2853) );
  AOI22X1 U859 ( .A0(n18183), .A1(\RAM<10><22> ), .B0(n18176), .B1(
        \RAM<8><22> ), .Y(n2837) );
  AOI22X1 U860 ( .A0(n18239), .A1(\RAM<2><22> ), .B0(n18232), .B1(\RAM<0><22> ), .Y(n2833) );
  AOI22X1 U861 ( .A0(n18183), .A1(\RAM<58><22> ), .B0(n18176), .B1(
        \RAM<56><22> ), .Y(n2847) );
  AOI22X1 U862 ( .A0(n18239), .A1(\RAM<50><22> ), .B0(n18232), .B1(
        \RAM<48><22> ), .Y(n2843) );
  AOI22X1 U863 ( .A0(n18183), .A1(\RAM<26><22> ), .B0(n18176), .B1(
        \RAM<24><22> ), .Y(n2867) );
  AOI22X1 U864 ( .A0(n18239), .A1(\RAM<18><22> ), .B0(n18232), .B1(
        \RAM<16><22> ), .Y(n2863) );
  AOI22X1 U865 ( .A0(n18182), .A1(\RAM<42><23> ), .B0(n18177), .B1(
        \RAM<40><23> ), .Y(n2813) );
  AOI22X1 U866 ( .A0(n18239), .A1(\RAM<34><23> ), .B0(n18233), .B1(
        \RAM<32><23> ), .Y(n2809) );
  AOI22X1 U867 ( .A0(n2079), .A1(\RAM<10><23> ), .B0(n18177), .B1(\RAM<8><23> ), .Y(n2793) );
  AOI22X1 U868 ( .A0(n2067), .A1(\RAM<2><23> ), .B0(n18233), .B1(\RAM<0><23> ), 
        .Y(n2789) );
  AOI22X1 U869 ( .A0(n2079), .A1(\RAM<58><23> ), .B0(n18177), .B1(
        \RAM<56><23> ), .Y(n2803) );
  AOI22X1 U870 ( .A0(n18240), .A1(\RAM<50><23> ), .B0(n18233), .B1(
        \RAM<48><23> ), .Y(n2799) );
  AOI22X1 U871 ( .A0(n18182), .A1(\RAM<26><23> ), .B0(n18177), .B1(
        \RAM<24><23> ), .Y(n2823) );
  AOI22X1 U872 ( .A0(n18241), .A1(\RAM<18><23> ), .B0(n18233), .B1(
        \RAM<16><23> ), .Y(n2819) );
  AOI22X1 U873 ( .A0(n18185), .A1(\RAM<42><24> ), .B0(n18177), .B1(
        \RAM<40><24> ), .Y(n2769) );
  AOI22X1 U874 ( .A0(n18240), .A1(\RAM<34><24> ), .B0(n18233), .B1(
        \RAM<32><24> ), .Y(n2765) );
  AOI22X1 U875 ( .A0(n2079), .A1(\RAM<10><24> ), .B0(n18177), .B1(\RAM<8><24> ), .Y(n2749) );
  AOI22X1 U876 ( .A0(n18241), .A1(\RAM<2><24> ), .B0(n18233), .B1(\RAM<0><24> ), .Y(n2745) );
  AOI22X1 U877 ( .A0(n18185), .A1(\RAM<58><24> ), .B0(n18177), .B1(
        \RAM<56><24> ), .Y(n2759) );
  AOI22X1 U878 ( .A0(n18241), .A1(\RAM<50><24> ), .B0(n18233), .B1(
        \RAM<48><24> ), .Y(n2755) );
  AOI22X1 U879 ( .A0(n18182), .A1(\RAM<26><24> ), .B0(n18177), .B1(
        \RAM<24><24> ), .Y(n2779) );
  AOI22X1 U880 ( .A0(n18239), .A1(\RAM<18><24> ), .B0(n18233), .B1(
        \RAM<16><24> ), .Y(n2775) );
  AOI22X1 U881 ( .A0(n18183), .A1(\RAM<42><25> ), .B0(n18177), .B1(
        \RAM<40><25> ), .Y(n2725) );
  AOI22X1 U882 ( .A0(n18241), .A1(\RAM<34><25> ), .B0(n18233), .B1(
        \RAM<32><25> ), .Y(n2721) );
  AOI22X1 U883 ( .A0(n2079), .A1(\RAM<10><25> ), .B0(n18177), .B1(\RAM<8><25> ), .Y(n2705) );
  AOI22X1 U884 ( .A0(n18239), .A1(\RAM<2><25> ), .B0(n18233), .B1(\RAM<0><25> ), .Y(n2701) );
  AOI22X1 U885 ( .A0(n18183), .A1(\RAM<58><25> ), .B0(n18177), .B1(
        \RAM<56><25> ), .Y(n2715) );
  AOI22X1 U886 ( .A0(n18241), .A1(\RAM<50><25> ), .B0(n18233), .B1(
        \RAM<48><25> ), .Y(n2711) );
  AOI22X1 U887 ( .A0(n18182), .A1(\RAM<26><25> ), .B0(n18177), .B1(
        \RAM<24><25> ), .Y(n2735) );
  AOI22X1 U888 ( .A0(n18240), .A1(\RAM<18><25> ), .B0(n18233), .B1(
        \RAM<16><25> ), .Y(n2731) );
  AOI22X1 U889 ( .A0(n18184), .A1(\RAM<10><26> ), .B0(n18174), .B1(
        \RAM<8><26> ), .Y(n2661) );
  AOI22X1 U890 ( .A0(n18240), .A1(\RAM<2><26> ), .B0(n18235), .B1(\RAM<0><26> ), .Y(n2657) );
  AOI22X1 U891 ( .A0(n18184), .A1(\RAM<42><26> ), .B0(n18174), .B1(
        \RAM<40><26> ), .Y(n2681) );
  AOI22X1 U892 ( .A0(n18240), .A1(\RAM<34><26> ), .B0(n18231), .B1(
        \RAM<32><26> ), .Y(n2677) );
  AOI22X1 U893 ( .A0(n18184), .A1(\RAM<58><26> ), .B0(n18174), .B1(
        \RAM<56><26> ), .Y(n2671) );
  AOI22X1 U894 ( .A0(n18240), .A1(\RAM<50><26> ), .B0(n18230), .B1(
        \RAM<48><26> ), .Y(n2667) );
  AOI22X1 U895 ( .A0(n18184), .A1(\RAM<26><26> ), .B0(n18177), .B1(
        \RAM<24><26> ), .Y(n2691) );
  AOI22X1 U896 ( .A0(n18240), .A1(\RAM<18><26> ), .B0(n18235), .B1(
        \RAM<16><26> ), .Y(n2687) );
  AOI22X1 U897 ( .A0(n18184), .A1(\RAM<10><27> ), .B0(n18177), .B1(
        \RAM<8><27> ), .Y(n2617) );
  AOI22X1 U898 ( .A0(n18240), .A1(\RAM<2><27> ), .B0(n18231), .B1(\RAM<0><27> ), .Y(n2613) );
  AOI22X1 U899 ( .A0(n18184), .A1(\RAM<42><27> ), .B0(n18177), .B1(
        \RAM<40><27> ), .Y(n2637) );
  AOI22X1 U900 ( .A0(n18240), .A1(\RAM<34><27> ), .B0(n18230), .B1(
        \RAM<32><27> ), .Y(n2633) );
  AOI22X1 U901 ( .A0(n18184), .A1(\RAM<58><27> ), .B0(n18174), .B1(
        \RAM<56><27> ), .Y(n2627) );
  AOI22X1 U902 ( .A0(n18240), .A1(\RAM<50><27> ), .B0(n18235), .B1(
        \RAM<48><27> ), .Y(n2623) );
  AOI22X1 U903 ( .A0(n18184), .A1(\RAM<26><27> ), .B0(n18174), .B1(
        \RAM<24><27> ), .Y(n2647) );
  AOI22X1 U904 ( .A0(n18240), .A1(\RAM<18><27> ), .B0(n18231), .B1(
        \RAM<16><27> ), .Y(n2643) );
  AOI22X1 U905 ( .A0(n18184), .A1(\RAM<10><28> ), .B0(n18176), .B1(
        \RAM<8><28> ), .Y(n2573) );
  AOI22X1 U906 ( .A0(n18240), .A1(\RAM<2><28> ), .B0(n2068), .B1(\RAM<0><28> ), 
        .Y(n2569) );
  AOI22X1 U907 ( .A0(n18184), .A1(\RAM<58><28> ), .B0(n18177), .B1(
        \RAM<56><28> ), .Y(n2583) );
  AOI22X1 U908 ( .A0(n18240), .A1(\RAM<50><28> ), .B0(n18230), .B1(
        \RAM<48><28> ), .Y(n2579) );
  AOI22X1 U909 ( .A0(n18184), .A1(\RAM<42><28> ), .B0(n18175), .B1(
        \RAM<40><28> ), .Y(n2593) );
  AOI22X1 U910 ( .A0(n18240), .A1(\RAM<34><28> ), .B0(n18231), .B1(
        \RAM<32><28> ), .Y(n2589) );
  AOI22X1 U911 ( .A0(n18184), .A1(\RAM<26><28> ), .B0(n18175), .B1(
        \RAM<24><28> ), .Y(n2603) );
  AOI22X1 U912 ( .A0(n18240), .A1(\RAM<18><28> ), .B0(n18235), .B1(
        \RAM<16><28> ), .Y(n2599) );
  AOI22X1 U913 ( .A0(n18185), .A1(\RAM<10><29> ), .B0(n18175), .B1(
        \RAM<8><29> ), .Y(n2529) );
  AOI22X1 U914 ( .A0(n2067), .A1(\RAM<2><29> ), .B0(n18234), .B1(\RAM<0><29> ), 
        .Y(n2525) );
  AOI22X1 U915 ( .A0(n18184), .A1(\RAM<58><29> ), .B0(n18175), .B1(
        \RAM<56><29> ), .Y(n2539) );
  AOI22X1 U916 ( .A0(n2067), .A1(\RAM<50><29> ), .B0(n18234), .B1(
        \RAM<48><29> ), .Y(n2535) );
  AOI22X1 U917 ( .A0(n18181), .A1(\RAM<42><29> ), .B0(n18174), .B1(
        \RAM<40><29> ), .Y(n2549) );
  AOI22X1 U918 ( .A0(n18239), .A1(\RAM<34><29> ), .B0(n18234), .B1(
        \RAM<32><29> ), .Y(n2545) );
  AOI22X1 U919 ( .A0(n18181), .A1(\RAM<26><29> ), .B0(n18174), .B1(
        \RAM<24><29> ), .Y(n2559) );
  AOI22X1 U920 ( .A0(n18239), .A1(\RAM<18><29> ), .B0(n18234), .B1(
        \RAM<16><29> ), .Y(n2555) );
  AOI22X1 U921 ( .A0(n18181), .A1(\RAM<10><30> ), .B0(n18174), .B1(
        \RAM<8><30> ), .Y(n2441) );
  AOI22X1 U922 ( .A0(n2067), .A1(\RAM<2><30> ), .B0(n18234), .B1(\RAM<0><30> ), 
        .Y(n2437) );
  AOI22X1 U923 ( .A0(n18184), .A1(\RAM<42><30> ), .B0(n18177), .B1(
        \RAM<40><30> ), .Y(n2461) );
  AOI22X1 U924 ( .A0(n18240), .A1(\RAM<34><30> ), .B0(n18234), .B1(
        \RAM<32><30> ), .Y(n2457) );
  AOI22X1 U925 ( .A0(n18184), .A1(\RAM<58><30> ), .B0(n18177), .B1(
        \RAM<56><30> ), .Y(n2451) );
  AOI22X1 U926 ( .A0(n18240), .A1(\RAM<50><30> ), .B0(n18234), .B1(
        \RAM<48><30> ), .Y(n2447) );
  AOI22X1 U927 ( .A0(n18186), .A1(\RAM<26><30> ), .B0(n18175), .B1(
        \RAM<24><30> ), .Y(n2471) );
  AOI22X1 U928 ( .A0(n18240), .A1(\RAM<18><30> ), .B0(n18234), .B1(
        \RAM<16><30> ), .Y(n2467) );
  AOI22X1 U929 ( .A0(n18185), .A1(\RAM<42><31> ), .B0(n18178), .B1(
        \RAM<40><31> ), .Y(n2417) );
  AOI22X1 U930 ( .A0(n18241), .A1(\RAM<34><31> ), .B0(n18233), .B1(
        \RAM<32><31> ), .Y(n2413) );
  AOI22X1 U931 ( .A0(n18185), .A1(\RAM<10><31> ), .B0(n18178), .B1(
        \RAM<8><31> ), .Y(n2397) );
  AOI22X1 U932 ( .A0(n18241), .A1(\RAM<2><31> ), .B0(n18233), .B1(\RAM<0><31> ), .Y(n2393) );
  AOI22X1 U933 ( .A0(n18185), .A1(\RAM<58><31> ), .B0(n18178), .B1(
        \RAM<56><31> ), .Y(n2407) );
  AOI22X1 U934 ( .A0(n18241), .A1(\RAM<50><31> ), .B0(n18233), .B1(
        \RAM<48><31> ), .Y(n2403) );
  AOI22X1 U935 ( .A0(n18185), .A1(\RAM<26><31> ), .B0(n18178), .B1(
        \RAM<24><31> ), .Y(n2427) );
  AOI22X1 U936 ( .A0(n18241), .A1(\RAM<18><31> ), .B0(n18233), .B1(
        \RAM<16><31> ), .Y(n2423) );
  AOI22X1 U937 ( .A0(n18182), .A1(\RAM<42><0> ), .B0(n18179), .B1(\RAM<40><0> ), .Y(n3473) );
  AOI22X1 U938 ( .A0(n18239), .A1(\RAM<34><0> ), .B0(n18233), .B1(\RAM<32><0> ), .Y(n3469) );
  AOI22X1 U939 ( .A0(n18184), .A1(\RAM<10><0> ), .B0(n2080), .B1(\RAM<8><0> ), 
        .Y(n3453) );
  AOI22X1 U940 ( .A0(n2067), .A1(\RAM<2><0> ), .B0(n18234), .B1(\RAM<0><0> ), 
        .Y(n3449) );
  AOI22X1 U941 ( .A0(n18185), .A1(\RAM<58><0> ), .B0(n18176), .B1(\RAM<56><0> ), .Y(n3463) );
  AOI22X1 U942 ( .A0(n18242), .A1(\RAM<50><0> ), .B0(n18234), .B1(\RAM<48><0> ), .Y(n3459) );
  AOI22X1 U943 ( .A0(n18185), .A1(\RAM<26><0> ), .B0(n18179), .B1(\RAM<24><0> ), .Y(n3489) );
  AOI22X1 U944 ( .A0(n18238), .A1(\RAM<18><0> ), .B0(n18233), .B1(\RAM<16><0> ), .Y(n3479) );
  AOI22X1 U945 ( .A0(n18181), .A1(\RAM<42><1> ), .B0(n18179), .B1(\RAM<40><1> ), .Y(n2989) );
  AOI22X1 U946 ( .A0(n18238), .A1(\RAM<34><1> ), .B0(n18235), .B1(\RAM<32><1> ), .Y(n2985) );
  AOI22X1 U947 ( .A0(n18186), .A1(\RAM<10><1> ), .B0(n18175), .B1(\RAM<8><1> ), 
        .Y(n2969) );
  AOI22X1 U948 ( .A0(n18238), .A1(\RAM<2><1> ), .B0(n18230), .B1(\RAM<0><1> ), 
        .Y(n2965) );
  AOI22X1 U949 ( .A0(n18181), .A1(\RAM<58><1> ), .B0(n18178), .B1(\RAM<56><1> ), .Y(n2979) );
  AOI22X1 U950 ( .A0(n18238), .A1(\RAM<50><1> ), .B0(n18231), .B1(\RAM<48><1> ), .Y(n2975) );
  AOI22X1 U951 ( .A0(n18184), .A1(\RAM<26><1> ), .B0(n18176), .B1(\RAM<24><1> ), .Y(n2999) );
  AOI22X1 U952 ( .A0(n18238), .A1(\RAM<18><1> ), .B0(n18230), .B1(\RAM<16><1> ), .Y(n2995) );
  AOI22X1 U953 ( .A0(n18167), .A1(\RAM<45><2> ), .B0(n18165), .B1(\RAM<41><2> ), .Y(n2504) );
  AOI22X1 U954 ( .A0(n18228), .A1(\RAM<37><2> ), .B0(n18220), .B1(\RAM<33><2> ), .Y(n2500) );
  AOI22X1 U955 ( .A0(n18171), .A1(\RAM<45><3> ), .B0(n18164), .B1(\RAM<41><3> ), .Y(n2372) );
  AOI22X1 U956 ( .A0(n18223), .A1(\RAM<37><3> ), .B0(n18218), .B1(\RAM<33><3> ), .Y(n2368) );
  AOI22X1 U957 ( .A0(n18170), .A1(\RAM<45><4> ), .B0(n18161), .B1(\RAM<41><4> ), .Y(n2328) );
  AOI22X1 U958 ( .A0(n18224), .A1(\RAM<37><4> ), .B0(n18220), .B1(\RAM<33><4> ), .Y(n2324) );
  AOI22X1 U959 ( .A0(n18172), .A1(\RAM<45><5> ), .B0(n18165), .B1(\RAM<41><5> ), .Y(n2284) );
  AOI22X1 U960 ( .A0(n18228), .A1(\RAM<37><5> ), .B0(n18221), .B1(\RAM<33><5> ), .Y(n2280) );
  AOI22X1 U961 ( .A0(n18172), .A1(\RAM<45><6> ), .B0(n18165), .B1(\RAM<41><6> ), .Y(n2240) );
  AOI22X1 U962 ( .A0(n18228), .A1(\RAM<37><6> ), .B0(n18221), .B1(\RAM<33><6> ), .Y(n2236) );
  AOI22X1 U963 ( .A0(n18172), .A1(\RAM<45><7> ), .B0(n18165), .B1(\RAM<41><7> ), .Y(n2196) );
  AOI22X1 U964 ( .A0(n18228), .A1(\RAM<37><7> ), .B0(n18221), .B1(\RAM<33><7> ), .Y(n2192) );
  AOI22X1 U965 ( .A0(n18170), .A1(\RAM<45><8> ), .B0(n18163), .B1(\RAM<41><8> ), .Y(n2152) );
  AOI22X1 U966 ( .A0(n18226), .A1(\RAM<37><8> ), .B0(n18220), .B1(\RAM<33><8> ), .Y(n2148) );
  AOI22X1 U967 ( .A0(n18168), .A1(\RAM<45><9> ), .B0(n18163), .B1(\RAM<41><9> ), .Y(n2107) );
  AOI22X1 U968 ( .A0(n18228), .A1(\RAM<37><9> ), .B0(n18221), .B1(\RAM<33><9> ), .Y(n2103) );
  AOI22X1 U969 ( .A0(n18167), .A1(\RAM<45><10> ), .B0(n18162), .B1(
        \RAM<41><10> ), .Y(n3428) );
  AOI22X1 U970 ( .A0(n18227), .A1(\RAM<37><10> ), .B0(n18220), .B1(
        \RAM<33><10> ), .Y(n3424) );
  AOI22X1 U971 ( .A0(n18167), .A1(\RAM<45><11> ), .B0(n18165), .B1(
        \RAM<41><11> ), .Y(n3384) );
  AOI22X1 U972 ( .A0(n18226), .A1(\RAM<37><11> ), .B0(n18219), .B1(
        \RAM<33><11> ), .Y(n3380) );
  AOI22X1 U973 ( .A0(n18168), .A1(\RAM<13><12> ), .B0(n18160), .B1(
        \RAM<9><12> ), .Y(n3320) );
  AOI22X1 U974 ( .A0(n18223), .A1(\RAM<5><12> ), .B0(n18216), .B1(\RAM<1><12> ), .Y(n3316) );
  AOI22X1 U975 ( .A0(n18168), .A1(\RAM<13><13> ), .B0(n18160), .B1(
        \RAM<9><13> ), .Y(n3276) );
  AOI22X1 U976 ( .A0(n18223), .A1(\RAM<5><13> ), .B0(n18216), .B1(\RAM<1><13> ), .Y(n3272) );
  AOI22X1 U977 ( .A0(n18168), .A1(\RAM<13><14> ), .B0(n18160), .B1(
        \RAM<9><14> ), .Y(n3232) );
  AOI22X1 U978 ( .A0(n18223), .A1(\RAM<5><14> ), .B0(n18216), .B1(\RAM<1><14> ), .Y(n3228) );
  AOI22X1 U979 ( .A0(n18169), .A1(\RAM<13><15> ), .B0(n18161), .B1(
        \RAM<9><15> ), .Y(n3188) );
  AOI22X1 U980 ( .A0(n18224), .A1(\RAM<5><15> ), .B0(n18217), .B1(\RAM<1><15> ), .Y(n3184) );
  AOI22X1 U981 ( .A0(n18169), .A1(\RAM<45><16> ), .B0(n18161), .B1(
        \RAM<41><16> ), .Y(n3164) );
  AOI22X1 U982 ( .A0(n18224), .A1(\RAM<37><16> ), .B0(n18217), .B1(
        \RAM<33><16> ), .Y(n3160) );
  AOI22X1 U983 ( .A0(n18169), .A1(\RAM<45><17> ), .B0(n18161), .B1(
        \RAM<41><17> ), .Y(n3120) );
  AOI22X1 U984 ( .A0(n18224), .A1(\RAM<37><17> ), .B0(n18217), .B1(
        \RAM<33><17> ), .Y(n3116) );
  AOI22X1 U985 ( .A0(n18170), .A1(\RAM<45><18> ), .B0(n18161), .B1(
        \RAM<41><18> ), .Y(n3076) );
  AOI22X1 U986 ( .A0(n18225), .A1(\RAM<37><18> ), .B0(n18217), .B1(
        \RAM<33><18> ), .Y(n3072) );
  AOI22X1 U987 ( .A0(n18170), .A1(\RAM<45><19> ), .B0(n18160), .B1(
        \RAM<41><19> ), .Y(n3032) );
  AOI22X1 U988 ( .A0(n18224), .A1(\RAM<37><19> ), .B0(n18216), .B1(
        \RAM<33><19> ), .Y(n3028) );
  AOI22X1 U989 ( .A0(n18171), .A1(\RAM<13><20> ), .B0(n18162), .B1(
        \RAM<9><20> ), .Y(n2924) );
  AOI22X1 U990 ( .A0(n18225), .A1(\RAM<5><20> ), .B0(n18218), .B1(\RAM<1><20> ), .Y(n2920) );
  AOI22X1 U991 ( .A0(n18171), .A1(\RAM<45><21> ), .B0(n18162), .B1(
        \RAM<41><21> ), .Y(n2900) );
  AOI22X1 U992 ( .A0(n18225), .A1(\RAM<37><21> ), .B0(n18218), .B1(
        \RAM<33><21> ), .Y(n2896) );
  AOI22X1 U993 ( .A0(n18171), .A1(\RAM<45><22> ), .B0(n18162), .B1(
        \RAM<41><22> ), .Y(n2856) );
  AOI22X1 U994 ( .A0(n18225), .A1(\RAM<37><22> ), .B0(n18218), .B1(
        \RAM<33><22> ), .Y(n2852) );
  AOI22X1 U995 ( .A0(n2081), .A1(\RAM<45><23> ), .B0(n18163), .B1(
        \RAM<41><23> ), .Y(n2812) );
  AOI22X1 U996 ( .A0(n18226), .A1(\RAM<37><23> ), .B0(n18219), .B1(
        \RAM<33><23> ), .Y(n2808) );
  AOI22X1 U997 ( .A0(n2081), .A1(\RAM<45><24> ), .B0(n18163), .B1(
        \RAM<41><24> ), .Y(n2768) );
  AOI22X1 U998 ( .A0(n18226), .A1(\RAM<37><24> ), .B0(n18219), .B1(
        \RAM<33><24> ), .Y(n2764) );
  AOI22X1 U999 ( .A0(n2081), .A1(\RAM<45><25> ), .B0(n18163), .B1(
        \RAM<41><25> ), .Y(n2724) );
  AOI22X1 U1000 ( .A0(n18226), .A1(\RAM<37><25> ), .B0(n18219), .B1(
        \RAM<33><25> ), .Y(n2720) );
  AOI22X1 U1001 ( .A0(n2081), .A1(\RAM<13><26> ), .B0(n18164), .B1(
        \RAM<9><26> ), .Y(n2660) );
  AOI22X1 U1002 ( .A0(n18227), .A1(\RAM<5><26> ), .B0(n18221), .B1(
        \RAM<1><26> ), .Y(n2656) );
  AOI22X1 U1003 ( .A0(n2081), .A1(\RAM<13><27> ), .B0(n18164), .B1(
        \RAM<9><27> ), .Y(n2616) );
  AOI22X1 U1004 ( .A0(n18227), .A1(\RAM<5><27> ), .B0(n18217), .B1(
        \RAM<1><27> ), .Y(n2612) );
  AOI22X1 U1005 ( .A0(n2081), .A1(\RAM<13><28> ), .B0(n18164), .B1(
        \RAM<9><28> ), .Y(n2572) );
  AOI22X1 U1006 ( .A0(n18227), .A1(\RAM<5><28> ), .B0(n2070), .B1(\RAM<1><28> ), .Y(n2568) );
  AOI22X1 U1007 ( .A0(n18172), .A1(\RAM<13><29> ), .B0(n18160), .B1(
        \RAM<9><29> ), .Y(n2528) );
  AOI22X1 U1008 ( .A0(n2069), .A1(\RAM<5><29> ), .B0(n18220), .B1(\RAM<1><29> ), .Y(n2524) );
  AOI22X1 U1009 ( .A0(n18169), .A1(\RAM<13><30> ), .B0(n18164), .B1(
        \RAM<9><30> ), .Y(n2440) );
  AOI22X1 U1010 ( .A0(n2069), .A1(\RAM<5><30> ), .B0(n18220), .B1(\RAM<1><30> ), .Y(n2436) );
  AOI22X1 U1011 ( .A0(n18169), .A1(\RAM<45><31> ), .B0(n18160), .B1(
        \RAM<41><31> ), .Y(n2416) );
  AOI22X1 U1012 ( .A0(n18223), .A1(\RAM<37><31> ), .B0(n18219), .B1(
        \RAM<33><31> ), .Y(n2412) );
  AOI22X1 U1013 ( .A0(n18167), .A1(\RAM<45><0> ), .B0(n18163), .B1(
        \RAM<41><0> ), .Y(n3472) );
  AOI22X1 U1014 ( .A0(n18227), .A1(\RAM<37><0> ), .B0(n18218), .B1(
        \RAM<33><0> ), .Y(n3468) );
  AOI22X1 U1015 ( .A0(n18170), .A1(\RAM<45><1> ), .B0(n18160), .B1(
        \RAM<41><1> ), .Y(n2988) );
  AOI22X1 U1016 ( .A0(n18224), .A1(\RAM<37><1> ), .B0(n18221), .B1(
        \RAM<33><1> ), .Y(n2984) );
  AOI22X1 U1017 ( .A0(n18153), .A1(\RAM<43><2> ), .B0(n18151), .B1(
        \RAM<46><2> ), .Y(n2503) );
  AOI22X1 U1018 ( .A0(n18213), .A1(\RAM<35><2> ), .B0(n18206), .B1(
        \RAM<38><2> ), .Y(n2499) );
  AOI22X1 U1019 ( .A0(n18157), .A1(\RAM<43><3> ), .B0(n18150), .B1(
        \RAM<46><3> ), .Y(n2371) );
  AOI22X1 U1020 ( .A0(n18212), .A1(\RAM<35><3> ), .B0(n18202), .B1(
        \RAM<38><3> ), .Y(n2367) );
  AOI22X1 U1021 ( .A0(n18156), .A1(\RAM<43><4> ), .B0(n18147), .B1(
        \RAM<46><4> ), .Y(n2327) );
  AOI22X1 U1022 ( .A0(n18209), .A1(\RAM<35><4> ), .B0(n18204), .B1(
        \RAM<38><4> ), .Y(n2323) );
  AOI22X1 U1023 ( .A0(n18158), .A1(\RAM<43><5> ), .B0(n18151), .B1(
        \RAM<46><5> ), .Y(n2283) );
  AOI22X1 U1024 ( .A0(n18210), .A1(\RAM<35><5> ), .B0(n18207), .B1(
        \RAM<38><5> ), .Y(n2279) );
  AOI22X1 U1025 ( .A0(n18158), .A1(\RAM<43><6> ), .B0(n18151), .B1(
        \RAM<46><6> ), .Y(n2239) );
  AOI22X1 U1026 ( .A0(n18214), .A1(\RAM<35><6> ), .B0(n18207), .B1(
        \RAM<38><6> ), .Y(n2235) );
  AOI22X1 U1027 ( .A0(n18158), .A1(\RAM<43><7> ), .B0(n18151), .B1(
        \RAM<46><7> ), .Y(n2195) );
  AOI22X1 U1028 ( .A0(n18211), .A1(\RAM<35><7> ), .B0(n18207), .B1(
        \RAM<38><7> ), .Y(n2191) );
  AOI22X1 U1029 ( .A0(n18156), .A1(\RAM<43><8> ), .B0(n18149), .B1(
        \RAM<46><8> ), .Y(n2151) );
  AOI22X1 U1030 ( .A0(n18209), .A1(\RAM<35><8> ), .B0(n18206), .B1(
        \RAM<38><8> ), .Y(n2147) );
  AOI22X1 U1031 ( .A0(n18154), .A1(\RAM<43><9> ), .B0(n18149), .B1(
        \RAM<46><9> ), .Y(n2106) );
  AOI22X1 U1032 ( .A0(n18211), .A1(\RAM<35><9> ), .B0(n18205), .B1(
        \RAM<38><9> ), .Y(n2102) );
  AOI22X1 U1033 ( .A0(n18153), .A1(\RAM<43><10> ), .B0(n18148), .B1(
        \RAM<46><10> ), .Y(n3427) );
  AOI22X1 U1034 ( .A0(n18209), .A1(\RAM<35><10> ), .B0(n18205), .B1(
        \RAM<38><10> ), .Y(n3423) );
  AOI22X1 U1035 ( .A0(n18153), .A1(\RAM<43><11> ), .B0(n18151), .B1(
        \RAM<46><11> ), .Y(n3383) );
  AOI22X1 U1036 ( .A0(n18209), .A1(\RAM<35><11> ), .B0(n18207), .B1(
        \RAM<38><11> ), .Y(n3379) );
  AOI22X1 U1037 ( .A0(n18154), .A1(\RAM<11><12> ), .B0(n18146), .B1(
        \RAM<14><12> ), .Y(n3319) );
  AOI22X1 U1038 ( .A0(n18210), .A1(\RAM<3><12> ), .B0(n18202), .B1(
        \RAM<6><12> ), .Y(n3315) );
  AOI22X1 U1039 ( .A0(n18154), .A1(\RAM<11><13> ), .B0(n18146), .B1(
        \RAM<14><13> ), .Y(n3275) );
  AOI22X1 U1040 ( .A0(n18210), .A1(\RAM<3><13> ), .B0(n18202), .B1(
        \RAM<6><13> ), .Y(n3271) );
  AOI22X1 U1041 ( .A0(n18154), .A1(\RAM<11><14> ), .B0(n18146), .B1(
        \RAM<14><14> ), .Y(n3231) );
  AOI22X1 U1042 ( .A0(n18210), .A1(\RAM<3><14> ), .B0(n18202), .B1(
        \RAM<6><14> ), .Y(n3227) );
  AOI22X1 U1043 ( .A0(n18155), .A1(\RAM<11><15> ), .B0(n18147), .B1(
        \RAM<14><15> ), .Y(n3187) );
  AOI22X1 U1044 ( .A0(n18211), .A1(\RAM<3><15> ), .B0(n18203), .B1(
        \RAM<6><15> ), .Y(n3183) );
  AOI22X1 U1045 ( .A0(n18155), .A1(\RAM<43><16> ), .B0(n18147), .B1(
        \RAM<46><16> ), .Y(n3163) );
  AOI22X1 U1046 ( .A0(n18211), .A1(\RAM<35><16> ), .B0(n18203), .B1(
        \RAM<38><16> ), .Y(n3159) );
  AOI22X1 U1047 ( .A0(n18155), .A1(\RAM<43><17> ), .B0(n18147), .B1(
        \RAM<46><17> ), .Y(n3119) );
  AOI22X1 U1048 ( .A0(n18211), .A1(\RAM<35><17> ), .B0(n18203), .B1(
        \RAM<38><17> ), .Y(n3115) );
  AOI22X1 U1049 ( .A0(n18156), .A1(\RAM<43><18> ), .B0(n18147), .B1(
        \RAM<46><18> ), .Y(n3075) );
  AOI22X1 U1050 ( .A0(n18211), .A1(\RAM<35><18> ), .B0(n18203), .B1(
        \RAM<38><18> ), .Y(n3071) );
  AOI22X1 U1051 ( .A0(n18156), .A1(\RAM<43><19> ), .B0(n18146), .B1(
        \RAM<46><19> ), .Y(n3031) );
  AOI22X1 U1052 ( .A0(n18210), .A1(\RAM<35><19> ), .B0(n18202), .B1(
        \RAM<38><19> ), .Y(n3027) );
  AOI22X1 U1053 ( .A0(n18157), .A1(\RAM<11><20> ), .B0(n18148), .B1(
        \RAM<14><20> ), .Y(n2923) );
  AOI22X1 U1054 ( .A0(n18212), .A1(\RAM<3><20> ), .B0(n18204), .B1(
        \RAM<6><20> ), .Y(n2919) );
  AOI22X1 U1055 ( .A0(n18157), .A1(\RAM<43><21> ), .B0(n18148), .B1(
        \RAM<46><21> ), .Y(n2899) );
  AOI22X1 U1056 ( .A0(n18212), .A1(\RAM<35><21> ), .B0(n18204), .B1(
        \RAM<38><21> ), .Y(n2895) );
  AOI22X1 U1057 ( .A0(n18157), .A1(\RAM<43><22> ), .B0(n18148), .B1(
        \RAM<46><22> ), .Y(n2855) );
  AOI22X1 U1058 ( .A0(n18212), .A1(\RAM<35><22> ), .B0(n18204), .B1(
        \RAM<38><22> ), .Y(n2851) );
  AOI22X1 U1059 ( .A0(n18154), .A1(\RAM<43><23> ), .B0(n18149), .B1(
        \RAM<46><23> ), .Y(n2811) );
  AOI22X1 U1060 ( .A0(n18213), .A1(\RAM<35><23> ), .B0(n18205), .B1(
        \RAM<38><23> ), .Y(n2807) );
  AOI22X1 U1061 ( .A0(n18156), .A1(\RAM<43><24> ), .B0(n18149), .B1(
        \RAM<46><24> ), .Y(n2767) );
  AOI22X1 U1062 ( .A0(n18213), .A1(\RAM<35><24> ), .B0(n18205), .B1(
        \RAM<38><24> ), .Y(n2763) );
  AOI22X1 U1063 ( .A0(n2083), .A1(\RAM<43><25> ), .B0(n18149), .B1(
        \RAM<46><25> ), .Y(n2723) );
  AOI22X1 U1064 ( .A0(n18213), .A1(\RAM<35><25> ), .B0(n18205), .B1(
        \RAM<38><25> ), .Y(n2719) );
  AOI22X1 U1065 ( .A0(n2083), .A1(\RAM<11><26> ), .B0(n18150), .B1(
        \RAM<14><26> ), .Y(n2659) );
  AOI22X1 U1066 ( .A0(n18214), .A1(\RAM<3><26> ), .B0(n18204), .B1(
        \RAM<6><26> ), .Y(n2655) );
  AOI22X1 U1067 ( .A0(n2083), .A1(\RAM<11><27> ), .B0(n18150), .B1(
        \RAM<14><27> ), .Y(n2615) );
  AOI22X1 U1068 ( .A0(n18214), .A1(\RAM<3><27> ), .B0(n18202), .B1(
        \RAM<6><27> ), .Y(n2611) );
  AOI22X1 U1069 ( .A0(n2083), .A1(\RAM<11><28> ), .B0(n18150), .B1(
        \RAM<14><28> ), .Y(n2571) );
  AOI22X1 U1070 ( .A0(n18214), .A1(\RAM<3><28> ), .B0(n18203), .B1(
        \RAM<6><28> ), .Y(n2567) );
  AOI22X1 U1071 ( .A0(n18158), .A1(\RAM<11><29> ), .B0(n18146), .B1(
        \RAM<14><29> ), .Y(n2527) );
  AOI22X1 U1072 ( .A0(n2071), .A1(\RAM<3><29> ), .B0(n18206), .B1(\RAM<6><29> ), .Y(n2523) );
  AOI22X1 U1073 ( .A0(n18156), .A1(\RAM<11><30> ), .B0(n18150), .B1(
        \RAM<14><30> ), .Y(n2439) );
  AOI22X1 U1074 ( .A0(n2071), .A1(\RAM<3><30> ), .B0(n18206), .B1(\RAM<6><30> ), .Y(n2435) );
  AOI22X1 U1075 ( .A0(n18155), .A1(\RAM<43><31> ), .B0(n18146), .B1(
        \RAM<46><31> ), .Y(n2415) );
  AOI22X1 U1076 ( .A0(n18213), .A1(\RAM<35><31> ), .B0(n18203), .B1(
        \RAM<38><31> ), .Y(n2411) );
  AOI22X1 U1077 ( .A0(n18153), .A1(\RAM<43><0> ), .B0(n18149), .B1(
        \RAM<46><0> ), .Y(n3471) );
  AOI22X1 U1078 ( .A0(n18209), .A1(\RAM<35><0> ), .B0(n18206), .B1(
        \RAM<38><0> ), .Y(n3467) );
  AOI22X1 U1079 ( .A0(n18156), .A1(\RAM<43><1> ), .B0(n18146), .B1(
        \RAM<46><1> ), .Y(n2987) );
  AOI22X1 U1080 ( .A0(n18214), .A1(\RAM<35><1> ), .B0(n18202), .B1(
        \RAM<38><1> ), .Y(n2983) );
  AOI22X1 U1081 ( .A0(n18142), .A1(\RAM<47><2> ), .B0(n18135), .B1(
        \RAM<44><2> ), .Y(n2502) );
  AOI22X1 U1082 ( .A0(n18141), .A1(\RAM<47><3> ), .B0(n18133), .B1(
        \RAM<44><3> ), .Y(n2370) );
  AOI22X1 U1083 ( .A0(n18141), .A1(\RAM<47><4> ), .B0(n18132), .B1(
        \RAM<44><4> ), .Y(n2326) );
  AOI22X1 U1084 ( .A0(n18144), .A1(\RAM<47><5> ), .B0(n18137), .B1(
        \RAM<44><5> ), .Y(n2282) );
  AOI22X1 U1085 ( .A0(n18144), .A1(\RAM<47><6> ), .B0(n18137), .B1(
        \RAM<44><6> ), .Y(n2238) );
  AOI22X1 U1086 ( .A0(n18144), .A1(\RAM<47><7> ), .B0(n18137), .B1(
        \RAM<44><7> ), .Y(n2194) );
  AOI22X1 U1087 ( .A0(n18139), .A1(\RAM<47><8> ), .B0(n18135), .B1(
        \RAM<44><8> ), .Y(n2150) );
  AOI22X1 U1088 ( .A0(n18144), .A1(\RAM<47><9> ), .B0(n18135), .B1(
        \RAM<44><9> ), .Y(n2105) );
  AOI22X1 U1089 ( .A0(n18139), .A1(\RAM<47><10> ), .B0(n18134), .B1(
        \RAM<44><10> ), .Y(n3426) );
  AOI22X1 U1090 ( .A0(n18139), .A1(\RAM<47><11> ), .B0(n18137), .B1(
        \RAM<44><11> ), .Y(n3382) );
  AOI22X1 U1091 ( .A0(n2085), .A1(\RAM<15><12> ), .B0(n18132), .B1(
        \RAM<12><12> ), .Y(n3318) );
  AOI22X1 U1092 ( .A0(n2085), .A1(\RAM<15><13> ), .B0(n18132), .B1(
        \RAM<12><13> ), .Y(n3274) );
  AOI22X1 U1093 ( .A0(n2085), .A1(\RAM<15><14> ), .B0(n18132), .B1(
        \RAM<12><14> ), .Y(n3230) );
  AOI22X1 U1094 ( .A0(n18140), .A1(\RAM<15><15> ), .B0(n18133), .B1(
        \RAM<12><15> ), .Y(n3186) );
  AOI22X1 U1095 ( .A0(n18140), .A1(\RAM<47><16> ), .B0(n18133), .B1(
        \RAM<44><16> ), .Y(n3162) );
  AOI22X1 U1096 ( .A0(n18140), .A1(\RAM<47><17> ), .B0(n18133), .B1(
        \RAM<44><17> ), .Y(n3118) );
  AOI22X1 U1097 ( .A0(n18143), .A1(\RAM<47><18> ), .B0(n18133), .B1(
        \RAM<44><18> ), .Y(n3074) );
  AOI22X1 U1098 ( .A0(n18143), .A1(\RAM<47><19> ), .B0(n18132), .B1(
        \RAM<44><19> ), .Y(n3030) );
  AOI22X1 U1099 ( .A0(n18141), .A1(\RAM<15><20> ), .B0(n18134), .B1(
        \RAM<12><20> ), .Y(n2922) );
  AOI22X1 U1100 ( .A0(n18141), .A1(\RAM<47><21> ), .B0(n18134), .B1(
        \RAM<44><21> ), .Y(n2898) );
  AOI22X1 U1101 ( .A0(n18141), .A1(\RAM<47><22> ), .B0(n18134), .B1(
        \RAM<44><22> ), .Y(n2854) );
  AOI22X1 U1102 ( .A0(n18142), .A1(\RAM<47><23> ), .B0(n18135), .B1(
        \RAM<44><23> ), .Y(n2810) );
  AOI22X1 U1103 ( .A0(n18142), .A1(\RAM<47><24> ), .B0(n18135), .B1(
        \RAM<44><24> ), .Y(n2766) );
  AOI22X1 U1104 ( .A0(n18142), .A1(\RAM<47><25> ), .B0(n18135), .B1(
        \RAM<44><25> ), .Y(n2722) );
  AOI22X1 U1105 ( .A0(n18143), .A1(\RAM<15><26> ), .B0(n18136), .B1(
        \RAM<12><26> ), .Y(n2658) );
  AOI22X1 U1106 ( .A0(n18143), .A1(\RAM<15><27> ), .B0(n18136), .B1(
        \RAM<12><27> ), .Y(n2614) );
  AOI22X1 U1107 ( .A0(n18143), .A1(\RAM<15><28> ), .B0(n18136), .B1(
        \RAM<12><28> ), .Y(n2570) );
  AOI22X1 U1108 ( .A0(n18142), .A1(\RAM<15><29> ), .B0(n18132), .B1(
        \RAM<12><29> ), .Y(n2526) );
  AOI22X1 U1109 ( .A0(n18142), .A1(\RAM<15><30> ), .B0(n18137), .B1(
        \RAM<12><30> ), .Y(n2438) );
  AOI22X1 U1110 ( .A0(n18144), .A1(\RAM<47><31> ), .B0(n18136), .B1(
        \RAM<44><31> ), .Y(n2414) );
  AOI22X1 U1111 ( .A0(n18139), .A1(\RAM<47><0> ), .B0(n18135), .B1(
        \RAM<44><0> ), .Y(n3470) );
  AOI22X1 U1112 ( .A0(n18142), .A1(\RAM<47><1> ), .B0(n18133), .B1(
        \RAM<44><1> ), .Y(n2986) );
  OAI21XL U1113 ( .A0(n3312), .A1(n3313), .B0(n18244), .Y(n3311) );
  NAND4X1 U1114 ( .A(n3314), .B(n3315), .C(n3316), .D(n3317), .Y(n3313) );
  NAND4X1 U1115 ( .A(n3318), .B(n3319), .C(n3320), .D(n3321), .Y(n3312) );
  AOI22X1 U1116 ( .A0(n18195), .A1(\RAM<7><12> ), .B0(n18189), .B1(
        \RAM<4><12> ), .Y(n3314) );
  OAI21XL U1117 ( .A0(n3268), .A1(n3269), .B0(n18244), .Y(n3267) );
  NAND4X1 U1118 ( .A(n3270), .B(n3271), .C(n3272), .D(n3273), .Y(n3269) );
  NAND4X1 U1119 ( .A(n3274), .B(n3275), .C(n3276), .D(n3277), .Y(n3268) );
  AOI22X1 U1120 ( .A0(n18195), .A1(\RAM<7><13> ), .B0(n18189), .B1(
        \RAM<4><13> ), .Y(n3270) );
  OAI21XL U1121 ( .A0(n3224), .A1(n3225), .B0(n18244), .Y(n3223) );
  NAND4X1 U1122 ( .A(n3226), .B(n3227), .C(n3228), .D(n3229), .Y(n3225) );
  NAND4X1 U1123 ( .A(n3230), .B(n3231), .C(n3232), .D(n3233), .Y(n3224) );
  AOI22X1 U1124 ( .A0(n18195), .A1(\RAM<7><14> ), .B0(n18189), .B1(
        \RAM<4><14> ), .Y(n3226) );
  OAI21XL U1125 ( .A0(n3180), .A1(n3181), .B0(n18244), .Y(n3179) );
  NAND4X1 U1126 ( .A(n3182), .B(n3183), .C(n3184), .D(n3185), .Y(n3181) );
  NAND4X1 U1127 ( .A(n3186), .B(n3187), .C(n3188), .D(n3189), .Y(n3180) );
  AOI22X1 U1128 ( .A0(n18196), .A1(\RAM<7><15> ), .B0(n18190), .B1(
        \RAM<4><15> ), .Y(n3182) );
  OAI21XL U1129 ( .A0(n2916), .A1(n2917), .B0(n18245), .Y(n2915) );
  NAND4X1 U1130 ( .A(n2918), .B(n2919), .C(n2920), .D(n2921), .Y(n2917) );
  NAND4X1 U1131 ( .A(n2922), .B(n2923), .C(n2924), .D(n2925), .Y(n2916) );
  AOI22X1 U1132 ( .A0(n18197), .A1(\RAM<7><20> ), .B0(n18189), .B1(
        \RAM<4><20> ), .Y(n2918) );
  OAI21XL U1133 ( .A0(n2652), .A1(n2653), .B0(n18245), .Y(n2651) );
  NAND4X1 U1134 ( .A(n2654), .B(n2655), .C(n2656), .D(n2657), .Y(n2653) );
  NAND4X1 U1135 ( .A(n2658), .B(n2659), .C(n2660), .D(n2661), .Y(n2652) );
  AOI22X1 U1136 ( .A0(n18199), .A1(\RAM<7><26> ), .B0(n18192), .B1(
        \RAM<4><26> ), .Y(n2654) );
  OAI21XL U1137 ( .A0(n2608), .A1(n2609), .B0(n18245), .Y(n2607) );
  NAND4X1 U1138 ( .A(n2610), .B(n2611), .C(n2612), .D(n2613), .Y(n2609) );
  NAND4X1 U1139 ( .A(n2614), .B(n2615), .C(n2616), .D(n2617), .Y(n2608) );
  AOI22X1 U1140 ( .A0(n18199), .A1(\RAM<7><27> ), .B0(n18191), .B1(
        \RAM<4><27> ), .Y(n2610) );
  OAI21XL U1141 ( .A0(n2564), .A1(n2565), .B0(n18245), .Y(n2563) );
  NAND4X1 U1142 ( .A(n2566), .B(n2567), .C(n2568), .D(n2569), .Y(n2565) );
  NAND4X1 U1143 ( .A(n2570), .B(n2571), .C(n2572), .D(n2573), .Y(n2564) );
  AOI22X1 U1144 ( .A0(n18199), .A1(\RAM<7><28> ), .B0(n18188), .B1(
        \RAM<4><28> ), .Y(n2566) );
  OAI21XL U1145 ( .A0(n2520), .A1(n2521), .B0(n18245), .Y(n2519) );
  NAND4X1 U1146 ( .A(n2522), .B(n2523), .C(n2524), .D(n2525), .Y(n2521) );
  NAND4X1 U1147 ( .A(n2526), .B(n2527), .C(n2528), .D(n2529), .Y(n2520) );
  AOI22X1 U1148 ( .A0(n18198), .A1(\RAM<7><29> ), .B0(n18191), .B1(
        \RAM<4><29> ), .Y(n2522) );
  OAI21XL U1149 ( .A0(n2432), .A1(n2433), .B0(n18245), .Y(n2431) );
  NAND4X1 U1150 ( .A(n2434), .B(n2435), .C(n2436), .D(n2437), .Y(n2433) );
  NAND4X1 U1151 ( .A(n2438), .B(n2439), .C(n2440), .D(n2441), .Y(n2432) );
  AOI22X1 U1152 ( .A0(n18197), .A1(\RAM<7><30> ), .B0(n18193), .B1(
        \RAM<4><30> ), .Y(n2434) );
  OAI21XL U1153 ( .A0(n2496), .A1(n2497), .B0(n18129), .Y(n2473) );
  NAND4X1 U1154 ( .A(n2498), .B(n2499), .C(n2500), .D(n2501), .Y(n2497) );
  NAND4X1 U1155 ( .A(n2502), .B(n2503), .C(n2504), .D(n2505), .Y(n2496) );
  AOI22X1 U1156 ( .A0(n18199), .A1(\RAM<39><2> ), .B0(n2074), .B1(\RAM<36><2> ), .Y(n2498) );
  OAI21XL U1157 ( .A0(n2364), .A1(n2365), .B0(n18129), .Y(n2341) );
  NAND4X1 U1158 ( .A(n2366), .B(n2367), .C(n2368), .D(n2369), .Y(n2365) );
  NAND4X1 U1159 ( .A(n2370), .B(n2371), .C(n2372), .D(n2373), .Y(n2364) );
  AOI22X1 U1160 ( .A0(n18196), .A1(\RAM<39><3> ), .B0(n18192), .B1(
        \RAM<36><3> ), .Y(n2366) );
  OAI21XL U1161 ( .A0(n2320), .A1(n2321), .B0(n18129), .Y(n2297) );
  NAND4X1 U1162 ( .A(n2322), .B(n2323), .C(n2324), .D(n2325), .Y(n2321) );
  NAND4X1 U1163 ( .A(n2326), .B(n2327), .C(n2328), .D(n2329), .Y(n2320) );
  AOI22X1 U1164 ( .A0(n18196), .A1(\RAM<39><4> ), .B0(n18192), .B1(
        \RAM<36><4> ), .Y(n2322) );
  OAI21XL U1165 ( .A0(n2276), .A1(n2277), .B0(n18129), .Y(n2253) );
  NAND4X1 U1166 ( .A(n2278), .B(n2279), .C(n2280), .D(n2281), .Y(n2277) );
  NAND4X1 U1167 ( .A(n2282), .B(n2283), .C(n2284), .D(n2285), .Y(n2276) );
  AOI22X1 U1168 ( .A0(n18200), .A1(\RAM<39><5> ), .B0(n18193), .B1(
        \RAM<36><5> ), .Y(n2278) );
  OAI21XL U1169 ( .A0(n2232), .A1(n2233), .B0(n18129), .Y(n2209) );
  NAND4X1 U1170 ( .A(n2234), .B(n2235), .C(n2236), .D(n2237), .Y(n2233) );
  NAND4X1 U1171 ( .A(n2238), .B(n2239), .C(n2240), .D(n2241), .Y(n2232) );
  AOI22X1 U1172 ( .A0(n18200), .A1(\RAM<39><6> ), .B0(n18193), .B1(
        \RAM<36><6> ), .Y(n2234) );
  OAI21XL U1173 ( .A0(n2188), .A1(n2189), .B0(n18129), .Y(n2165) );
  NAND4X1 U1174 ( .A(n2190), .B(n2191), .C(n2192), .D(n2193), .Y(n2189) );
  NAND4X1 U1175 ( .A(n2194), .B(n2195), .C(n2196), .D(n2197), .Y(n2188) );
  AOI22X1 U1176 ( .A0(n18200), .A1(\RAM<39><7> ), .B0(n18193), .B1(
        \RAM<36><7> ), .Y(n2190) );
  OAI21XL U1177 ( .A0(n2144), .A1(n2145), .B0(n18129), .Y(n2121) );
  NAND4X1 U1178 ( .A(n2146), .B(n2147), .C(n2148), .D(n2149), .Y(n2145) );
  NAND4X1 U1179 ( .A(n2150), .B(n2151), .C(n2152), .D(n2153), .Y(n2144) );
  AOI22X1 U1180 ( .A0(n18200), .A1(\RAM<39><8> ), .B0(n18188), .B1(
        \RAM<36><8> ), .Y(n2146) );
  OAI21XL U1181 ( .A0(n2098), .A1(n2099), .B0(n18129), .Y(n2057) );
  NAND4X1 U1182 ( .A(n2101), .B(n2102), .C(n2103), .D(n2104), .Y(n2099) );
  NAND4X1 U1183 ( .A(n2105), .B(n2106), .C(n2107), .D(n2108), .Y(n2098) );
  AOI22X1 U1184 ( .A0(n18199), .A1(\RAM<39><9> ), .B0(n18193), .B1(
        \RAM<36><9> ), .Y(n2101) );
  OAI21XL U1185 ( .A0(n3420), .A1(n3421), .B0(n18128), .Y(n3397) );
  NAND4X1 U1186 ( .A(n3422), .B(n3423), .C(n3424), .D(n3425), .Y(n3421) );
  NAND4X1 U1187 ( .A(n3426), .B(n3427), .C(n3428), .D(n3429), .Y(n3420) );
  AOI22X1 U1188 ( .A0(n18198), .A1(\RAM<39><10> ), .B0(n18188), .B1(
        \RAM<36><10> ), .Y(n3422) );
  OAI21XL U1189 ( .A0(n3376), .A1(n3377), .B0(n18128), .Y(n3353) );
  NAND4X1 U1190 ( .A(n3378), .B(n3379), .C(n3380), .D(n3381), .Y(n3377) );
  NAND4X1 U1191 ( .A(n3382), .B(n3383), .C(n3384), .D(n3385), .Y(n3376) );
  AOI22X1 U1192 ( .A0(n18197), .A1(\RAM<39><11> ), .B0(n18188), .B1(
        \RAM<36><11> ), .Y(n3378) );
  OAI21XL U1193 ( .A0(n3156), .A1(n3157), .B0(n18128), .Y(n3133) );
  NAND4X1 U1194 ( .A(n3158), .B(n3159), .C(n3160), .D(n3161), .Y(n3157) );
  NAND4X1 U1195 ( .A(n3162), .B(n3163), .C(n3164), .D(n3165), .Y(n3156) );
  AOI22X1 U1196 ( .A0(n18196), .A1(\RAM<39><16> ), .B0(n18190), .B1(
        \RAM<36><16> ), .Y(n3158) );
  OAI21XL U1197 ( .A0(n3112), .A1(n3113), .B0(n18128), .Y(n3089) );
  NAND4X1 U1198 ( .A(n3114), .B(n3115), .C(n3116), .D(n3117), .Y(n3113) );
  NAND4X1 U1199 ( .A(n3118), .B(n3119), .C(n3120), .D(n3121), .Y(n3112) );
  AOI22X1 U1200 ( .A0(n18196), .A1(\RAM<39><17> ), .B0(n18190), .B1(
        \RAM<36><17> ), .Y(n3114) );
  OAI21XL U1201 ( .A0(n3068), .A1(n3069), .B0(n18128), .Y(n3045) );
  NAND4X1 U1202 ( .A(n3070), .B(n3071), .C(n3072), .D(n3073), .Y(n3069) );
  NAND4X1 U1203 ( .A(n3074), .B(n3075), .C(n3076), .D(n3077), .Y(n3068) );
  AOI22X1 U1204 ( .A0(n18200), .A1(\RAM<39><18> ), .B0(n18190), .B1(
        \RAM<36><18> ), .Y(n3070) );
  OAI21XL U1205 ( .A0(n3024), .A1(n3025), .B0(n18128), .Y(n3001) );
  NAND4X1 U1206 ( .A(n3026), .B(n3027), .C(n3028), .D(n3029), .Y(n3025) );
  NAND4X1 U1207 ( .A(n3030), .B(n3031), .C(n3032), .D(n3033), .Y(n3024) );
  AOI22X1 U1208 ( .A0(n18196), .A1(\RAM<39><19> ), .B0(n18189), .B1(
        \RAM<36><19> ), .Y(n3026) );
  OAI21XL U1209 ( .A0(n2892), .A1(n2893), .B0(n18129), .Y(n2869) );
  NAND4X1 U1210 ( .A(n2894), .B(n2895), .C(n2896), .D(n2897), .Y(n2893) );
  NAND4X1 U1211 ( .A(n2898), .B(n2899), .C(n2900), .D(n2901), .Y(n2892) );
  AOI22X1 U1212 ( .A0(n18197), .A1(\RAM<39><21> ), .B0(n18189), .B1(
        \RAM<36><21> ), .Y(n2894) );
  OAI21XL U1213 ( .A0(n2848), .A1(n2849), .B0(n18129), .Y(n2825) );
  NAND4X1 U1214 ( .A(n2850), .B(n2851), .C(n2852), .D(n2853), .Y(n2849) );
  NAND4X1 U1215 ( .A(n2854), .B(n2855), .C(n2856), .D(n2857), .Y(n2848) );
  AOI22X1 U1216 ( .A0(n18197), .A1(\RAM<39><22> ), .B0(n18190), .B1(
        \RAM<36><22> ), .Y(n2850) );
  OAI21XL U1217 ( .A0(n2804), .A1(n2805), .B0(n18129), .Y(n2781) );
  NAND4X1 U1218 ( .A(n2806), .B(n2807), .C(n2808), .D(n2809), .Y(n2805) );
  NAND4X1 U1219 ( .A(n2810), .B(n2811), .C(n2812), .D(n2813), .Y(n2804) );
  AOI22X1 U1220 ( .A0(n18198), .A1(\RAM<39><23> ), .B0(n18191), .B1(
        \RAM<36><23> ), .Y(n2806) );
  OAI21XL U1221 ( .A0(n2760), .A1(n2761), .B0(n18129), .Y(n2737) );
  NAND4X1 U1222 ( .A(n2762), .B(n2763), .C(n2764), .D(n2765), .Y(n2761) );
  NAND4X1 U1223 ( .A(n2766), .B(n2767), .C(n2768), .D(n2769), .Y(n2760) );
  AOI22X1 U1224 ( .A0(n18198), .A1(\RAM<39><24> ), .B0(n18191), .B1(
        \RAM<36><24> ), .Y(n2762) );
  OAI21XL U1225 ( .A0(n2716), .A1(n2717), .B0(n18129), .Y(n2693) );
  NAND4X1 U1226 ( .A(n2718), .B(n2719), .C(n2720), .D(n2721), .Y(n2717) );
  NAND4X1 U1227 ( .A(n2722), .B(n2723), .C(n2724), .D(n2725), .Y(n2716) );
  AOI22X1 U1228 ( .A0(n18198), .A1(\RAM<39><25> ), .B0(n18191), .B1(
        \RAM<36><25> ), .Y(n2718) );
  OAI21XL U1229 ( .A0(n2408), .A1(n2409), .B0(n18129), .Y(n2385) );
  NAND4X1 U1230 ( .A(n2410), .B(n2411), .C(n2412), .D(n2413), .Y(n2409) );
  NAND4X1 U1231 ( .A(n2414), .B(n2415), .C(n2416), .D(n2417), .Y(n2408) );
  AOI22X1 U1232 ( .A0(n18195), .A1(\RAM<39><31> ), .B0(n18192), .B1(
        \RAM<36><31> ), .Y(n2410) );
  OAI21XL U1233 ( .A0(n3464), .A1(n3465), .B0(n18128), .Y(n3441) );
  NAND4X1 U1234 ( .A(n3466), .B(n3467), .C(n3468), .D(n3469), .Y(n3465) );
  NAND4X1 U1235 ( .A(n3470), .B(n3471), .C(n3472), .D(n3473), .Y(n3464) );
  AOI22X1 U1236 ( .A0(n18199), .A1(\RAM<39><0> ), .B0(n18188), .B1(
        \RAM<36><0> ), .Y(n3466) );
  OAI21XL U1237 ( .A0(n2980), .A1(n2981), .B0(n18129), .Y(n2957) );
  NAND4X1 U1238 ( .A(n2982), .B(n2983), .C(n2984), .D(n2985), .Y(n2981) );
  NAND4X1 U1239 ( .A(n2986), .B(n2987), .C(n2988), .D(n2989), .Y(n2980) );
  AOI22X1 U1240 ( .A0(n18195), .A1(\RAM<39><1> ), .B0(n2074), .B1(\RAM<36><1> ), .Y(n2982) );
  NAND4X1 U1241 ( .A(n2482), .B(n2483), .C(n2484), .D(n2485), .Y(n2476) );
  AOI22X1 U1242 ( .A0(n18140), .A1(\RAM<15><2> ), .B0(n18133), .B1(
        \RAM<12><2> ), .Y(n2482) );
  AOI22X1 U1243 ( .A0(n2083), .A1(\RAM<11><2> ), .B0(n18147), .B1(\RAM<14><2> ), .Y(n2483) );
  AOI22X1 U1244 ( .A0(n2081), .A1(\RAM<13><2> ), .B0(n18161), .B1(\RAM<9><2> ), 
        .Y(n2484) );
  NAND4X1 U1245 ( .A(n2492), .B(n2493), .C(n2494), .D(n2495), .Y(n2486) );
  AOI22X1 U1246 ( .A0(n18143), .A1(\RAM<63><2> ), .B0(n18136), .B1(
        \RAM<60><2> ), .Y(n2492) );
  AOI22X1 U1247 ( .A0(n18158), .A1(\RAM<59><2> ), .B0(n18151), .B1(
        \RAM<62><2> ), .Y(n2493) );
  AOI22X1 U1248 ( .A0(n18172), .A1(\RAM<61><2> ), .B0(n18165), .B1(
        \RAM<57><2> ), .Y(n2494) );
  NAND4X1 U1249 ( .A(n2512), .B(n2513), .C(n2514), .D(n2515), .Y(n2506) );
  AOI22X1 U1250 ( .A0(n18140), .A1(\RAM<31><2> ), .B0(n18135), .B1(
        \RAM<28><2> ), .Y(n2512) );
  AOI22X1 U1251 ( .A0(n2083), .A1(\RAM<27><2> ), .B0(n18149), .B1(\RAM<30><2> ), .Y(n2513) );
  AOI22X1 U1252 ( .A0(n18169), .A1(\RAM<29><2> ), .B0(n18163), .B1(
        \RAM<25><2> ), .Y(n2514) );
  NAND4X1 U1253 ( .A(n2350), .B(n2351), .C(n2352), .D(n2353), .Y(n2344) );
  AOI22X1 U1254 ( .A0(n18144), .A1(\RAM<15><3> ), .B0(n18136), .B1(
        \RAM<12><3> ), .Y(n2350) );
  AOI22X1 U1255 ( .A0(n18155), .A1(\RAM<11><3> ), .B0(n18147), .B1(
        \RAM<14><3> ), .Y(n2351) );
  AOI22X1 U1256 ( .A0(n18169), .A1(\RAM<13><3> ), .B0(n18161), .B1(\RAM<9><3> ), .Y(n2352) );
  NAND4X1 U1257 ( .A(n2360), .B(n2361), .C(n2362), .D(n2363), .Y(n2354) );
  AOI22X1 U1258 ( .A0(n18139), .A1(\RAM<63><3> ), .B0(n18132), .B1(
        \RAM<60><3> ), .Y(n2360) );
  AOI22X1 U1259 ( .A0(n18154), .A1(\RAM<59><3> ), .B0(n18150), .B1(
        \RAM<62><3> ), .Y(n2361) );
  AOI22X1 U1260 ( .A0(n18168), .A1(\RAM<61><3> ), .B0(n18164), .B1(
        \RAM<57><3> ), .Y(n2362) );
  NAND4X1 U1261 ( .A(n2380), .B(n2381), .C(n2382), .D(n2383), .Y(n2374) );
  AOI22X1 U1262 ( .A0(n18141), .A1(\RAM<31><3> ), .B0(n18136), .B1(
        \RAM<28><3> ), .Y(n2380) );
  AOI22X1 U1263 ( .A0(n18156), .A1(\RAM<27><3> ), .B0(n18146), .B1(
        \RAM<30><3> ), .Y(n2381) );
  AOI22X1 U1264 ( .A0(n18170), .A1(\RAM<29><3> ), .B0(n18160), .B1(
        \RAM<25><3> ), .Y(n2382) );
  NAND4X1 U1265 ( .A(n2306), .B(n2307), .C(n2308), .D(n2309), .Y(n2300) );
  AOI22X1 U1266 ( .A0(n18139), .A1(\RAM<15><4> ), .B0(n18133), .B1(
        \RAM<12><4> ), .Y(n2306) );
  AOI22X1 U1267 ( .A0(n18154), .A1(\RAM<11><4> ), .B0(n18150), .B1(
        \RAM<14><4> ), .Y(n2307) );
  AOI22X1 U1268 ( .A0(n18168), .A1(\RAM<13><4> ), .B0(n18160), .B1(\RAM<9><4> ), .Y(n2308) );
  NAND4X1 U1269 ( .A(n2316), .B(n2317), .C(n2318), .D(n2319), .Y(n2310) );
  AOI22X1 U1270 ( .A0(n2085), .A1(\RAM<63><4> ), .B0(n18136), .B1(\RAM<60><4> ), .Y(n2316) );
  AOI22X1 U1271 ( .A0(n18157), .A1(\RAM<59><4> ), .B0(n18147), .B1(
        \RAM<62><4> ), .Y(n2317) );
  AOI22X1 U1272 ( .A0(n18171), .A1(\RAM<61><4> ), .B0(n18161), .B1(
        \RAM<57><4> ), .Y(n2318) );
  NAND4X1 U1273 ( .A(n2336), .B(n2337), .C(n2338), .D(n2339), .Y(n2330) );
  AOI22X1 U1274 ( .A0(n18144), .A1(\RAM<31><4> ), .B0(n18133), .B1(
        \RAM<28><4> ), .Y(n2336) );
  AOI22X1 U1275 ( .A0(n18155), .A1(\RAM<27><4> ), .B0(n18150), .B1(
        \RAM<30><4> ), .Y(n2337) );
  AOI22X1 U1276 ( .A0(n18169), .A1(\RAM<29><4> ), .B0(n18164), .B1(
        \RAM<25><4> ), .Y(n2338) );
  NAND4X1 U1277 ( .A(n2262), .B(n2263), .C(n2264), .D(n2265), .Y(n2256) );
  AOI22X1 U1278 ( .A0(n18144), .A1(\RAM<15><5> ), .B0(n18137), .B1(
        \RAM<12><5> ), .Y(n2262) );
  AOI22X1 U1279 ( .A0(n18158), .A1(\RAM<11><5> ), .B0(n18151), .B1(
        \RAM<14><5> ), .Y(n2263) );
  AOI22X1 U1280 ( .A0(n18172), .A1(\RAM<13><5> ), .B0(n18165), .B1(\RAM<9><5> ), .Y(n2264) );
  NAND4X1 U1281 ( .A(n2272), .B(n2273), .C(n2274), .D(n2275), .Y(n2266) );
  AOI22X1 U1282 ( .A0(n18144), .A1(\RAM<63><5> ), .B0(n18137), .B1(
        \RAM<60><5> ), .Y(n2272) );
  AOI22X1 U1283 ( .A0(n18158), .A1(\RAM<59><5> ), .B0(n18151), .B1(
        \RAM<62><5> ), .Y(n2273) );
  AOI22X1 U1284 ( .A0(n18172), .A1(\RAM<61><5> ), .B0(n18165), .B1(
        \RAM<57><5> ), .Y(n2274) );
  NAND4X1 U1285 ( .A(n2292), .B(n2293), .C(n2294), .D(n2295), .Y(n2286) );
  AOI22X1 U1286 ( .A0(n18144), .A1(\RAM<31><5> ), .B0(n18137), .B1(
        \RAM<28><5> ), .Y(n2292) );
  AOI22X1 U1287 ( .A0(n18158), .A1(\RAM<27><5> ), .B0(n18151), .B1(
        \RAM<30><5> ), .Y(n2293) );
  AOI22X1 U1288 ( .A0(n18172), .A1(\RAM<29><5> ), .B0(n18165), .B1(
        \RAM<25><5> ), .Y(n2294) );
  NAND4X1 U1289 ( .A(n2218), .B(n2219), .C(n2220), .D(n2221), .Y(n2212) );
  AOI22X1 U1290 ( .A0(n18144), .A1(\RAM<15><6> ), .B0(n18137), .B1(
        \RAM<12><6> ), .Y(n2218) );
  AOI22X1 U1291 ( .A0(n18158), .A1(\RAM<11><6> ), .B0(n18151), .B1(
        \RAM<14><6> ), .Y(n2219) );
  AOI22X1 U1292 ( .A0(n18172), .A1(\RAM<13><6> ), .B0(n18165), .B1(\RAM<9><6> ), .Y(n2220) );
  NAND4X1 U1293 ( .A(n2228), .B(n2229), .C(n2230), .D(n2231), .Y(n2222) );
  AOI22X1 U1294 ( .A0(n18144), .A1(\RAM<63><6> ), .B0(n18137), .B1(
        \RAM<60><6> ), .Y(n2228) );
  AOI22X1 U1295 ( .A0(n18158), .A1(\RAM<59><6> ), .B0(n18151), .B1(
        \RAM<62><6> ), .Y(n2229) );
  AOI22X1 U1296 ( .A0(n18172), .A1(\RAM<61><6> ), .B0(n18165), .B1(
        \RAM<57><6> ), .Y(n2230) );
  NAND4X1 U1297 ( .A(n2248), .B(n2249), .C(n2250), .D(n2251), .Y(n2242) );
  AOI22X1 U1298 ( .A0(n18144), .A1(\RAM<31><6> ), .B0(n18137), .B1(
        \RAM<28><6> ), .Y(n2248) );
  AOI22X1 U1299 ( .A0(n18158), .A1(\RAM<27><6> ), .B0(n18151), .B1(
        \RAM<30><6> ), .Y(n2249) );
  AOI22X1 U1300 ( .A0(n18172), .A1(\RAM<29><6> ), .B0(n18165), .B1(
        \RAM<25><6> ), .Y(n2250) );
  NAND4X1 U1301 ( .A(n2174), .B(n2175), .C(n2176), .D(n2177), .Y(n2168) );
  AOI22X1 U1302 ( .A0(n18144), .A1(\RAM<15><7> ), .B0(n18137), .B1(
        \RAM<12><7> ), .Y(n2174) );
  AOI22X1 U1303 ( .A0(n18158), .A1(\RAM<11><7> ), .B0(n18151), .B1(
        \RAM<14><7> ), .Y(n2175) );
  AOI22X1 U1304 ( .A0(n18172), .A1(\RAM<13><7> ), .B0(n18165), .B1(\RAM<9><7> ), .Y(n2176) );
  NAND4X1 U1305 ( .A(n2184), .B(n2185), .C(n2186), .D(n2187), .Y(n2178) );
  AOI22X1 U1306 ( .A0(n18144), .A1(\RAM<63><7> ), .B0(n18137), .B1(
        \RAM<60><7> ), .Y(n2184) );
  AOI22X1 U1307 ( .A0(n18158), .A1(\RAM<59><7> ), .B0(n18151), .B1(
        \RAM<62><7> ), .Y(n2185) );
  AOI22X1 U1308 ( .A0(n18172), .A1(\RAM<61><7> ), .B0(n18165), .B1(
        \RAM<57><7> ), .Y(n2186) );
  NAND4X1 U1309 ( .A(n2204), .B(n2205), .C(n2206), .D(n2207), .Y(n2198) );
  AOI22X1 U1310 ( .A0(n18144), .A1(\RAM<31><7> ), .B0(n18137), .B1(
        \RAM<28><7> ), .Y(n2204) );
  AOI22X1 U1311 ( .A0(n18158), .A1(\RAM<27><7> ), .B0(n18151), .B1(
        \RAM<30><7> ), .Y(n2205) );
  AOI22X1 U1312 ( .A0(n18172), .A1(\RAM<29><7> ), .B0(n18165), .B1(
        \RAM<25><7> ), .Y(n2206) );
  NAND4X1 U1313 ( .A(n3406), .B(n3407), .C(n3408), .D(n3409), .Y(n3400) );
  AOI22X1 U1314 ( .A0(n18139), .A1(\RAM<15><10> ), .B0(n18135), .B1(
        \RAM<12><10> ), .Y(n3406) );
  AOI22X1 U1315 ( .A0(n18153), .A1(\RAM<11><10> ), .B0(n18149), .B1(
        \RAM<14><10> ), .Y(n3407) );
  AOI22X1 U1316 ( .A0(n18167), .A1(\RAM<13><10> ), .B0(n18163), .B1(
        \RAM<9><10> ), .Y(n3408) );
  NAND4X1 U1317 ( .A(n3416), .B(n3417), .C(n3418), .D(n3419), .Y(n3410) );
  AOI22X1 U1318 ( .A0(n18139), .A1(\RAM<63><10> ), .B0(n18137), .B1(
        \RAM<60><10> ), .Y(n3416) );
  AOI22X1 U1319 ( .A0(n18153), .A1(\RAM<59><10> ), .B0(n18151), .B1(
        \RAM<62><10> ), .Y(n3417) );
  AOI22X1 U1320 ( .A0(n18167), .A1(\RAM<61><10> ), .B0(n18165), .B1(
        \RAM<57><10> ), .Y(n3418) );
  NAND4X1 U1321 ( .A(n3436), .B(n3437), .C(n3438), .D(n3439), .Y(n3430) );
  AOI22X1 U1322 ( .A0(n18139), .A1(\RAM<31><10> ), .B0(n18135), .B1(
        \RAM<28><10> ), .Y(n3436) );
  AOI22X1 U1323 ( .A0(n18153), .A1(\RAM<27><10> ), .B0(n18148), .B1(
        \RAM<30><10> ), .Y(n3437) );
  AOI22X1 U1324 ( .A0(n18167), .A1(\RAM<29><10> ), .B0(n18162), .B1(
        \RAM<25><10> ), .Y(n3438) );
  NAND4X1 U1325 ( .A(n3362), .B(n3363), .C(n3364), .D(n3365), .Y(n3356) );
  AOI22X1 U1326 ( .A0(n18139), .A1(\RAM<15><11> ), .B0(n18134), .B1(
        \RAM<12><11> ), .Y(n3362) );
  AOI22X1 U1327 ( .A0(n18153), .A1(\RAM<11><11> ), .B0(n18148), .B1(
        \RAM<14><11> ), .Y(n3363) );
  AOI22X1 U1328 ( .A0(n18167), .A1(\RAM<13><11> ), .B0(n18162), .B1(
        \RAM<9><11> ), .Y(n3364) );
  NAND4X1 U1329 ( .A(n3372), .B(n3373), .C(n3374), .D(n3375), .Y(n3366) );
  AOI22X1 U1330 ( .A0(n18139), .A1(\RAM<63><11> ), .B0(n18135), .B1(
        \RAM<60><11> ), .Y(n3372) );
  AOI22X1 U1331 ( .A0(n18153), .A1(\RAM<59><11> ), .B0(n18149), .B1(
        \RAM<62><11> ), .Y(n3373) );
  AOI22X1 U1332 ( .A0(n18167), .A1(\RAM<61><11> ), .B0(n18163), .B1(
        \RAM<57><11> ), .Y(n3374) );
  NAND4X1 U1333 ( .A(n3392), .B(n3393), .C(n3394), .D(n3395), .Y(n3386) );
  AOI22X1 U1334 ( .A0(n18139), .A1(\RAM<31><11> ), .B0(n18134), .B1(
        \RAM<28><11> ), .Y(n3392) );
  AOI22X1 U1335 ( .A0(n18153), .A1(\RAM<27><11> ), .B0(n18149), .B1(
        \RAM<30><11> ), .Y(n3393) );
  AOI22X1 U1336 ( .A0(n18167), .A1(\RAM<29><11> ), .B0(n18163), .B1(
        \RAM<25><11> ), .Y(n3394) );
  NAND4X1 U1337 ( .A(n3338), .B(n3339), .C(n3340), .D(n3341), .Y(n3332) );
  AOI22X1 U1338 ( .A0(n18141), .A1(\RAM<47><12> ), .B0(n18132), .B1(
        \RAM<44><12> ), .Y(n3338) );
  AOI22X1 U1339 ( .A0(n18154), .A1(\RAM<43><12> ), .B0(n18146), .B1(
        \RAM<46><12> ), .Y(n3339) );
  AOI22X1 U1340 ( .A0(n18168), .A1(\RAM<45><12> ), .B0(n18160), .B1(
        \RAM<41><12> ), .Y(n3340) );
  NAND4X1 U1341 ( .A(n3328), .B(n3329), .C(n3330), .D(n3331), .Y(n3322) );
  AOI22X1 U1342 ( .A0(n18139), .A1(\RAM<63><12> ), .B0(n18132), .B1(
        \RAM<60><12> ), .Y(n3328) );
  AOI22X1 U1343 ( .A0(n18154), .A1(\RAM<59><12> ), .B0(n18146), .B1(
        \RAM<62><12> ), .Y(n3329) );
  AOI22X1 U1344 ( .A0(n18168), .A1(\RAM<61><12> ), .B0(n18160), .B1(
        \RAM<57><12> ), .Y(n3330) );
  NAND4X1 U1345 ( .A(n3348), .B(n3349), .C(n3350), .D(n3351), .Y(n3342) );
  AOI22X1 U1346 ( .A0(n18141), .A1(\RAM<31><12> ), .B0(n18132), .B1(
        \RAM<28><12> ), .Y(n3348) );
  AOI22X1 U1347 ( .A0(n18154), .A1(\RAM<27><12> ), .B0(n18146), .B1(
        \RAM<30><12> ), .Y(n3349) );
  AOI22X1 U1348 ( .A0(n18168), .A1(\RAM<29><12> ), .B0(n18160), .B1(
        \RAM<25><12> ), .Y(n3350) );
  NAND4X1 U1349 ( .A(n3294), .B(n3295), .C(n3296), .D(n3297), .Y(n3288) );
  AOI22X1 U1350 ( .A0(n18144), .A1(\RAM<47><13> ), .B0(n18132), .B1(
        \RAM<44><13> ), .Y(n3294) );
  AOI22X1 U1351 ( .A0(n18154), .A1(\RAM<43><13> ), .B0(n18146), .B1(
        \RAM<46><13> ), .Y(n3295) );
  AOI22X1 U1352 ( .A0(n18168), .A1(\RAM<45><13> ), .B0(n18160), .B1(
        \RAM<41><13> ), .Y(n3296) );
  NAND4X1 U1353 ( .A(n3284), .B(n3285), .C(n3286), .D(n3287), .Y(n3278) );
  AOI22X1 U1354 ( .A0(n2085), .A1(\RAM<63><13> ), .B0(n18132), .B1(
        \RAM<60><13> ), .Y(n3284) );
  AOI22X1 U1355 ( .A0(n18154), .A1(\RAM<59><13> ), .B0(n18146), .B1(
        \RAM<62><13> ), .Y(n3285) );
  AOI22X1 U1356 ( .A0(n18168), .A1(\RAM<61><13> ), .B0(n18160), .B1(
        \RAM<57><13> ), .Y(n3286) );
  NAND4X1 U1357 ( .A(n3304), .B(n3305), .C(n3306), .D(n3307), .Y(n3298) );
  AOI22X1 U1358 ( .A0(n18144), .A1(\RAM<31><13> ), .B0(n18132), .B1(
        \RAM<28><13> ), .Y(n3304) );
  AOI22X1 U1359 ( .A0(n18154), .A1(\RAM<27><13> ), .B0(n18146), .B1(
        \RAM<30><13> ), .Y(n3305) );
  AOI22X1 U1360 ( .A0(n18168), .A1(\RAM<29><13> ), .B0(n18160), .B1(
        \RAM<25><13> ), .Y(n3306) );
  NAND4X1 U1361 ( .A(n3250), .B(n3251), .C(n3252), .D(n3253), .Y(n3244) );
  AOI22X1 U1362 ( .A0(n18139), .A1(\RAM<47><14> ), .B0(n18132), .B1(
        \RAM<44><14> ), .Y(n3250) );
  AOI22X1 U1363 ( .A0(n18154), .A1(\RAM<43><14> ), .B0(n18146), .B1(
        \RAM<46><14> ), .Y(n3251) );
  AOI22X1 U1364 ( .A0(n18168), .A1(\RAM<45><14> ), .B0(n18160), .B1(
        \RAM<41><14> ), .Y(n3252) );
  NAND4X1 U1365 ( .A(n3240), .B(n3241), .C(n3242), .D(n3243), .Y(n3234) );
  AOI22X1 U1366 ( .A0(n2085), .A1(\RAM<63><14> ), .B0(n18132), .B1(
        \RAM<60><14> ), .Y(n3240) );
  AOI22X1 U1367 ( .A0(n18154), .A1(\RAM<59><14> ), .B0(n18146), .B1(
        \RAM<62><14> ), .Y(n3241) );
  AOI22X1 U1368 ( .A0(n18168), .A1(\RAM<61><14> ), .B0(n18160), .B1(
        \RAM<57><14> ), .Y(n3242) );
  NAND4X1 U1369 ( .A(n3260), .B(n3261), .C(n3262), .D(n3263), .Y(n3254) );
  AOI22X1 U1370 ( .A0(n18139), .A1(\RAM<31><14> ), .B0(n18132), .B1(
        \RAM<28><14> ), .Y(n3260) );
  AOI22X1 U1371 ( .A0(n18154), .A1(\RAM<27><14> ), .B0(n18146), .B1(
        \RAM<30><14> ), .Y(n3261) );
  AOI22X1 U1372 ( .A0(n18168), .A1(\RAM<29><14> ), .B0(n18160), .B1(
        \RAM<25><14> ), .Y(n3262) );
  NAND4X1 U1373 ( .A(n3206), .B(n3207), .C(n3208), .D(n3209), .Y(n3200) );
  AOI22X1 U1374 ( .A0(n18140), .A1(\RAM<47><15> ), .B0(n18133), .B1(
        \RAM<44><15> ), .Y(n3206) );
  AOI22X1 U1375 ( .A0(n18155), .A1(\RAM<43><15> ), .B0(n18147), .B1(
        \RAM<46><15> ), .Y(n3207) );
  AOI22X1 U1376 ( .A0(n18169), .A1(\RAM<45><15> ), .B0(n18161), .B1(
        \RAM<41><15> ), .Y(n3208) );
  NAND4X1 U1377 ( .A(n3196), .B(n3197), .C(n3198), .D(n3199), .Y(n3190) );
  AOI22X1 U1378 ( .A0(n18140), .A1(\RAM<63><15> ), .B0(n18133), .B1(
        \RAM<60><15> ), .Y(n3196) );
  AOI22X1 U1379 ( .A0(n18155), .A1(\RAM<59><15> ), .B0(n18147), .B1(
        \RAM<62><15> ), .Y(n3197) );
  AOI22X1 U1380 ( .A0(n18169), .A1(\RAM<61><15> ), .B0(n18161), .B1(
        \RAM<57><15> ), .Y(n3198) );
  NAND4X1 U1381 ( .A(n3216), .B(n3217), .C(n3218), .D(n3219), .Y(n3210) );
  AOI22X1 U1382 ( .A0(n18140), .A1(\RAM<31><15> ), .B0(n18133), .B1(
        \RAM<28><15> ), .Y(n3216) );
  AOI22X1 U1383 ( .A0(n18155), .A1(\RAM<27><15> ), .B0(n18147), .B1(
        \RAM<30><15> ), .Y(n3217) );
  AOI22X1 U1384 ( .A0(n18169), .A1(\RAM<29><15> ), .B0(n18161), .B1(
        \RAM<25><15> ), .Y(n3218) );
  NAND4X1 U1385 ( .A(n3142), .B(n3143), .C(n3144), .D(n3145), .Y(n3136) );
  AOI22X1 U1386 ( .A0(n18140), .A1(\RAM<15><16> ), .B0(n18133), .B1(
        \RAM<12><16> ), .Y(n3142) );
  AOI22X1 U1387 ( .A0(n18155), .A1(\RAM<11><16> ), .B0(n18147), .B1(
        \RAM<14><16> ), .Y(n3143) );
  AOI22X1 U1388 ( .A0(n18169), .A1(\RAM<13><16> ), .B0(n18161), .B1(
        \RAM<9><16> ), .Y(n3144) );
  NAND4X1 U1389 ( .A(n3152), .B(n3153), .C(n3154), .D(n3155), .Y(n3146) );
  AOI22X1 U1390 ( .A0(n18140), .A1(\RAM<63><16> ), .B0(n18133), .B1(
        \RAM<60><16> ), .Y(n3152) );
  AOI22X1 U1391 ( .A0(n18155), .A1(\RAM<59><16> ), .B0(n18147), .B1(
        \RAM<62><16> ), .Y(n3153) );
  AOI22X1 U1392 ( .A0(n18169), .A1(\RAM<61><16> ), .B0(n18161), .B1(
        \RAM<57><16> ), .Y(n3154) );
  NAND4X1 U1393 ( .A(n3172), .B(n3173), .C(n3174), .D(n3175), .Y(n3166) );
  AOI22X1 U1394 ( .A0(n18140), .A1(\RAM<31><16> ), .B0(n18133), .B1(
        \RAM<28><16> ), .Y(n3172) );
  AOI22X1 U1395 ( .A0(n18155), .A1(\RAM<27><16> ), .B0(n18147), .B1(
        \RAM<30><16> ), .Y(n3173) );
  AOI22X1 U1396 ( .A0(n18169), .A1(\RAM<29><16> ), .B0(n18161), .B1(
        \RAM<25><16> ), .Y(n3174) );
  NAND4X1 U1397 ( .A(n3098), .B(n3099), .C(n3100), .D(n3101), .Y(n3092) );
  AOI22X1 U1398 ( .A0(n18140), .A1(\RAM<15><17> ), .B0(n18133), .B1(
        \RAM<12><17> ), .Y(n3098) );
  AOI22X1 U1399 ( .A0(n18155), .A1(\RAM<11><17> ), .B0(n18147), .B1(
        \RAM<14><17> ), .Y(n3099) );
  AOI22X1 U1400 ( .A0(n18169), .A1(\RAM<13><17> ), .B0(n18161), .B1(
        \RAM<9><17> ), .Y(n3100) );
  NAND4X1 U1401 ( .A(n3108), .B(n3109), .C(n3110), .D(n3111), .Y(n3102) );
  AOI22X1 U1402 ( .A0(n18140), .A1(\RAM<63><17> ), .B0(n18133), .B1(
        \RAM<60><17> ), .Y(n3108) );
  AOI22X1 U1403 ( .A0(n18155), .A1(\RAM<59><17> ), .B0(n18147), .B1(
        \RAM<62><17> ), .Y(n3109) );
  AOI22X1 U1404 ( .A0(n18169), .A1(\RAM<61><17> ), .B0(n18161), .B1(
        \RAM<57><17> ), .Y(n3110) );
  NAND4X1 U1405 ( .A(n3128), .B(n3129), .C(n3130), .D(n3131), .Y(n3122) );
  AOI22X1 U1406 ( .A0(n18140), .A1(\RAM<31><17> ), .B0(n18133), .B1(
        \RAM<28><17> ), .Y(n3128) );
  AOI22X1 U1407 ( .A0(n18155), .A1(\RAM<27><17> ), .B0(n18147), .B1(
        \RAM<30><17> ), .Y(n3129) );
  AOI22X1 U1408 ( .A0(n18169), .A1(\RAM<29><17> ), .B0(n18161), .B1(
        \RAM<25><17> ), .Y(n3130) );
  NAND4X1 U1409 ( .A(n3054), .B(n3055), .C(n3056), .D(n3057), .Y(n3048) );
  AOI22X1 U1410 ( .A0(n18140), .A1(\RAM<15><18> ), .B0(n18136), .B1(
        \RAM<12><18> ), .Y(n3054) );
  AOI22X1 U1411 ( .A0(n18156), .A1(\RAM<11><18> ), .B0(n18150), .B1(
        \RAM<14><18> ), .Y(n3055) );
  AOI22X1 U1412 ( .A0(n18170), .A1(\RAM<13><18> ), .B0(n18164), .B1(
        \RAM<9><18> ), .Y(n3056) );
  NAND4X1 U1413 ( .A(n3064), .B(n3065), .C(n3066), .D(n3067), .Y(n3058) );
  AOI22X1 U1414 ( .A0(n18142), .A1(\RAM<63><18> ), .B0(n18132), .B1(
        \RAM<60><18> ), .Y(n3064) );
  AOI22X1 U1415 ( .A0(n18156), .A1(\RAM<59><18> ), .B0(n18146), .B1(
        \RAM<62><18> ), .Y(n3065) );
  AOI22X1 U1416 ( .A0(n18170), .A1(\RAM<61><18> ), .B0(n18160), .B1(
        \RAM<57><18> ), .Y(n3066) );
  NAND4X1 U1417 ( .A(n3084), .B(n3085), .C(n3086), .D(n3087), .Y(n3078) );
  AOI22X1 U1418 ( .A0(n18142), .A1(\RAM<31><18> ), .B0(n18133), .B1(
        \RAM<28><18> ), .Y(n3084) );
  AOI22X1 U1419 ( .A0(n18156), .A1(\RAM<27><18> ), .B0(n18147), .B1(
        \RAM<30><18> ), .Y(n3085) );
  AOI22X1 U1420 ( .A0(n18170), .A1(\RAM<29><18> ), .B0(n18161), .B1(
        \RAM<25><18> ), .Y(n3086) );
  NAND4X1 U1421 ( .A(n3010), .B(n3011), .C(n3012), .D(n3013), .Y(n3004) );
  AOI22X1 U1422 ( .A0(n18142), .A1(\RAM<15><19> ), .B0(n2086), .B1(
        \RAM<12><19> ), .Y(n3010) );
  AOI22X1 U1423 ( .A0(n18156), .A1(\RAM<11><19> ), .B0(n2084), .B1(
        \RAM<14><19> ), .Y(n3011) );
  AOI22X1 U1424 ( .A0(n18170), .A1(\RAM<13><19> ), .B0(n2082), .B1(
        \RAM<9><19> ), .Y(n3012) );
  NAND4X1 U1425 ( .A(n3020), .B(n3021), .C(n3022), .D(n3023), .Y(n3014) );
  AOI22X1 U1426 ( .A0(n18143), .A1(\RAM<63><19> ), .B0(n18133), .B1(
        \RAM<60><19> ), .Y(n3020) );
  AOI22X1 U1427 ( .A0(n18156), .A1(\RAM<59><19> ), .B0(n18147), .B1(
        \RAM<62><19> ), .Y(n3021) );
  AOI22X1 U1428 ( .A0(n18170), .A1(\RAM<61><19> ), .B0(n18161), .B1(
        \RAM<57><19> ), .Y(n3022) );
  NAND4X1 U1429 ( .A(n3040), .B(n3041), .C(n3042), .D(n3043), .Y(n3034) );
  AOI22X1 U1430 ( .A0(n18140), .A1(\RAM<31><19> ), .B0(n18132), .B1(
        \RAM<28><19> ), .Y(n3040) );
  AOI22X1 U1431 ( .A0(n18156), .A1(\RAM<27><19> ), .B0(n18146), .B1(
        \RAM<30><19> ), .Y(n3041) );
  AOI22X1 U1432 ( .A0(n18170), .A1(\RAM<29><19> ), .B0(n18160), .B1(
        \RAM<25><19> ), .Y(n3042) );
  NAND4X1 U1433 ( .A(n2942), .B(n2943), .C(n2944), .D(n2945), .Y(n2936) );
  AOI22X1 U1434 ( .A0(n18141), .A1(\RAM<47><20> ), .B0(n18134), .B1(
        \RAM<44><20> ), .Y(n2942) );
  AOI22X1 U1435 ( .A0(n18157), .A1(\RAM<43><20> ), .B0(n18148), .B1(
        \RAM<46><20> ), .Y(n2943) );
  AOI22X1 U1436 ( .A0(n18171), .A1(\RAM<45><20> ), .B0(n18162), .B1(
        \RAM<41><20> ), .Y(n2944) );
  NAND4X1 U1437 ( .A(n2932), .B(n2933), .C(n2934), .D(n2935), .Y(n2926) );
  AOI22X1 U1438 ( .A0(n18141), .A1(\RAM<63><20> ), .B0(n18134), .B1(
        \RAM<60><20> ), .Y(n2932) );
  AOI22X1 U1439 ( .A0(n18157), .A1(\RAM<59><20> ), .B0(n18148), .B1(
        \RAM<62><20> ), .Y(n2933) );
  AOI22X1 U1440 ( .A0(n18171), .A1(\RAM<61><20> ), .B0(n18162), .B1(
        \RAM<57><20> ), .Y(n2934) );
  NAND4X1 U1441 ( .A(n2952), .B(n2953), .C(n2954), .D(n2955), .Y(n2946) );
  AOI22X1 U1442 ( .A0(n18141), .A1(\RAM<31><20> ), .B0(n18134), .B1(
        \RAM<28><20> ), .Y(n2952) );
  AOI22X1 U1443 ( .A0(n18157), .A1(\RAM<27><20> ), .B0(n18148), .B1(
        \RAM<30><20> ), .Y(n2953) );
  AOI22X1 U1444 ( .A0(n18171), .A1(\RAM<29><20> ), .B0(n18162), .B1(
        \RAM<25><20> ), .Y(n2954) );
  NAND4X1 U1445 ( .A(n2878), .B(n2879), .C(n2880), .D(n2881), .Y(n2872) );
  AOI22X1 U1446 ( .A0(n18141), .A1(\RAM<15><21> ), .B0(n18134), .B1(
        \RAM<12><21> ), .Y(n2878) );
  AOI22X1 U1447 ( .A0(n18157), .A1(\RAM<11><21> ), .B0(n18148), .B1(
        \RAM<14><21> ), .Y(n2879) );
  AOI22X1 U1448 ( .A0(n18171), .A1(\RAM<13><21> ), .B0(n18162), .B1(
        \RAM<9><21> ), .Y(n2880) );
  NAND4X1 U1449 ( .A(n2888), .B(n2889), .C(n2890), .D(n2891), .Y(n2882) );
  AOI22X1 U1450 ( .A0(n18141), .A1(\RAM<63><21> ), .B0(n18134), .B1(
        \RAM<60><21> ), .Y(n2888) );
  AOI22X1 U1451 ( .A0(n18157), .A1(\RAM<59><21> ), .B0(n18148), .B1(
        \RAM<62><21> ), .Y(n2889) );
  AOI22X1 U1452 ( .A0(n18171), .A1(\RAM<61><21> ), .B0(n18162), .B1(
        \RAM<57><21> ), .Y(n2890) );
  NAND4X1 U1453 ( .A(n2908), .B(n2909), .C(n2910), .D(n2911), .Y(n2902) );
  AOI22X1 U1454 ( .A0(n18141), .A1(\RAM<31><21> ), .B0(n18134), .B1(
        \RAM<28><21> ), .Y(n2908) );
  AOI22X1 U1455 ( .A0(n18157), .A1(\RAM<27><21> ), .B0(n18148), .B1(
        \RAM<30><21> ), .Y(n2909) );
  AOI22X1 U1456 ( .A0(n18171), .A1(\RAM<29><21> ), .B0(n18162), .B1(
        \RAM<25><21> ), .Y(n2910) );
  NAND4X1 U1457 ( .A(n2834), .B(n2835), .C(n2836), .D(n2837), .Y(n2828) );
  AOI22X1 U1458 ( .A0(n18141), .A1(\RAM<15><22> ), .B0(n18134), .B1(
        \RAM<12><22> ), .Y(n2834) );
  AOI22X1 U1459 ( .A0(n18157), .A1(\RAM<11><22> ), .B0(n18148), .B1(
        \RAM<14><22> ), .Y(n2835) );
  AOI22X1 U1460 ( .A0(n18171), .A1(\RAM<13><22> ), .B0(n18162), .B1(
        \RAM<9><22> ), .Y(n2836) );
  NAND4X1 U1461 ( .A(n2844), .B(n2845), .C(n2846), .D(n2847), .Y(n2838) );
  AOI22X1 U1462 ( .A0(n18141), .A1(\RAM<63><22> ), .B0(n18134), .B1(
        \RAM<60><22> ), .Y(n2844) );
  AOI22X1 U1463 ( .A0(n18157), .A1(\RAM<59><22> ), .B0(n18148), .B1(
        \RAM<62><22> ), .Y(n2845) );
  AOI22X1 U1464 ( .A0(n18171), .A1(\RAM<61><22> ), .B0(n18162), .B1(
        \RAM<57><22> ), .Y(n2846) );
  NAND4X1 U1465 ( .A(n2864), .B(n2865), .C(n2866), .D(n2867), .Y(n2858) );
  AOI22X1 U1466 ( .A0(n18141), .A1(\RAM<31><22> ), .B0(n18134), .B1(
        \RAM<28><22> ), .Y(n2864) );
  AOI22X1 U1467 ( .A0(n18157), .A1(\RAM<27><22> ), .B0(n18148), .B1(
        \RAM<30><22> ), .Y(n2865) );
  AOI22X1 U1468 ( .A0(n18171), .A1(\RAM<29><22> ), .B0(n18162), .B1(
        \RAM<25><22> ), .Y(n2866) );
  NAND4X1 U1469 ( .A(n2790), .B(n2791), .C(n2792), .D(n2793), .Y(n2784) );
  AOI22X1 U1470 ( .A0(n18142), .A1(\RAM<15><23> ), .B0(n18135), .B1(
        \RAM<12><23> ), .Y(n2790) );
  AOI22X1 U1471 ( .A0(n18157), .A1(\RAM<11><23> ), .B0(n18149), .B1(
        \RAM<14><23> ), .Y(n2791) );
  AOI22X1 U1472 ( .A0(n18171), .A1(\RAM<13><23> ), .B0(n18163), .B1(
        \RAM<9><23> ), .Y(n2792) );
  NAND4X1 U1473 ( .A(n2800), .B(n2801), .C(n2802), .D(n2803), .Y(n2794) );
  AOI22X1 U1474 ( .A0(n18142), .A1(\RAM<63><23> ), .B0(n18135), .B1(
        \RAM<60><23> ), .Y(n2800) );
  AOI22X1 U1475 ( .A0(n18157), .A1(\RAM<59><23> ), .B0(n18149), .B1(
        \RAM<62><23> ), .Y(n2801) );
  AOI22X1 U1476 ( .A0(n18171), .A1(\RAM<61><23> ), .B0(n18163), .B1(
        \RAM<57><23> ), .Y(n2802) );
  NAND4X1 U1477 ( .A(n2820), .B(n2821), .C(n2822), .D(n2823), .Y(n2814) );
  AOI22X1 U1478 ( .A0(n18142), .A1(\RAM<31><23> ), .B0(n18135), .B1(
        \RAM<28><23> ), .Y(n2820) );
  AOI22X1 U1479 ( .A0(n2083), .A1(\RAM<27><23> ), .B0(n18149), .B1(
        \RAM<30><23> ), .Y(n2821) );
  AOI22X1 U1480 ( .A0(n18168), .A1(\RAM<29><23> ), .B0(n18163), .B1(
        \RAM<25><23> ), .Y(n2822) );
  NAND4X1 U1481 ( .A(n2746), .B(n2747), .C(n2748), .D(n2749), .Y(n2740) );
  AOI22X1 U1482 ( .A0(n18142), .A1(\RAM<15><24> ), .B0(n18135), .B1(
        \RAM<12><24> ), .Y(n2746) );
  AOI22X1 U1483 ( .A0(n18155), .A1(\RAM<11><24> ), .B0(n18149), .B1(
        \RAM<14><24> ), .Y(n2747) );
  AOI22X1 U1484 ( .A0(n18170), .A1(\RAM<13><24> ), .B0(n18163), .B1(
        \RAM<9><24> ), .Y(n2748) );
  NAND4X1 U1485 ( .A(n2756), .B(n2757), .C(n2758), .D(n2759), .Y(n2750) );
  AOI22X1 U1486 ( .A0(n18142), .A1(\RAM<63><24> ), .B0(n18135), .B1(
        \RAM<60><24> ), .Y(n2756) );
  AOI22X1 U1487 ( .A0(n18156), .A1(\RAM<59><24> ), .B0(n18149), .B1(
        \RAM<62><24> ), .Y(n2757) );
  AOI22X1 U1488 ( .A0(n18170), .A1(\RAM<61><24> ), .B0(n18163), .B1(
        \RAM<57><24> ), .Y(n2758) );
  NAND4X1 U1489 ( .A(n2776), .B(n2777), .C(n2778), .D(n2779), .Y(n2770) );
  AOI22X1 U1490 ( .A0(n18142), .A1(\RAM<31><24> ), .B0(n18135), .B1(
        \RAM<28><24> ), .Y(n2776) );
  AOI22X1 U1491 ( .A0(n2083), .A1(\RAM<27><24> ), .B0(n18149), .B1(
        \RAM<30><24> ), .Y(n2777) );
  AOI22X1 U1492 ( .A0(n18170), .A1(\RAM<29><24> ), .B0(n18163), .B1(
        \RAM<25><24> ), .Y(n2778) );
  NAND4X1 U1493 ( .A(n2702), .B(n2703), .C(n2704), .D(n2705), .Y(n2696) );
  AOI22X1 U1494 ( .A0(n18142), .A1(\RAM<15><25> ), .B0(n18135), .B1(
        \RAM<12><25> ), .Y(n2702) );
  AOI22X1 U1495 ( .A0(n18154), .A1(\RAM<11><25> ), .B0(n18149), .B1(
        \RAM<14><25> ), .Y(n2703) );
  AOI22X1 U1496 ( .A0(n18168), .A1(\RAM<13><25> ), .B0(n18163), .B1(
        \RAM<9><25> ), .Y(n2704) );
  NAND4X1 U1497 ( .A(n2712), .B(n2713), .C(n2714), .D(n2715), .Y(n2706) );
  AOI22X1 U1498 ( .A0(n18142), .A1(\RAM<63><25> ), .B0(n18135), .B1(
        \RAM<60><25> ), .Y(n2712) );
  AOI22X1 U1499 ( .A0(n18157), .A1(\RAM<59><25> ), .B0(n18149), .B1(
        \RAM<62><25> ), .Y(n2713) );
  AOI22X1 U1500 ( .A0(n18169), .A1(\RAM<61><25> ), .B0(n18163), .B1(
        \RAM<57><25> ), .Y(n2714) );
  NAND4X1 U1501 ( .A(n2732), .B(n2733), .C(n2734), .D(n2735), .Y(n2726) );
  AOI22X1 U1502 ( .A0(n18142), .A1(\RAM<31><25> ), .B0(n18135), .B1(
        \RAM<28><25> ), .Y(n2732) );
  AOI22X1 U1503 ( .A0(n2083), .A1(\RAM<27><25> ), .B0(n18149), .B1(
        \RAM<30><25> ), .Y(n2733) );
  AOI22X1 U1504 ( .A0(n2081), .A1(\RAM<29><25> ), .B0(n18163), .B1(
        \RAM<25><25> ), .Y(n2734) );
  NAND4X1 U1505 ( .A(n2678), .B(n2679), .C(n2680), .D(n2681), .Y(n2672) );
  AOI22X1 U1506 ( .A0(n18143), .A1(\RAM<47><26> ), .B0(n18136), .B1(
        \RAM<44><26> ), .Y(n2678) );
  AOI22X1 U1507 ( .A0(n18158), .A1(\RAM<43><26> ), .B0(n18150), .B1(
        \RAM<46><26> ), .Y(n2679) );
  AOI22X1 U1508 ( .A0(n18172), .A1(\RAM<45><26> ), .B0(n18164), .B1(
        \RAM<41><26> ), .Y(n2680) );
  NAND4X1 U1509 ( .A(n2668), .B(n2669), .C(n2670), .D(n2671), .Y(n2662) );
  AOI22X1 U1510 ( .A0(n18143), .A1(\RAM<63><26> ), .B0(n18136), .B1(
        \RAM<60><26> ), .Y(n2668) );
  AOI22X1 U1511 ( .A0(n18155), .A1(\RAM<59><26> ), .B0(n18150), .B1(
        \RAM<62><26> ), .Y(n2669) );
  AOI22X1 U1512 ( .A0(n18171), .A1(\RAM<61><26> ), .B0(n18164), .B1(
        \RAM<57><26> ), .Y(n2670) );
  NAND4X1 U1513 ( .A(n2688), .B(n2689), .C(n2690), .D(n2691), .Y(n2682) );
  AOI22X1 U1514 ( .A0(n18143), .A1(\RAM<31><26> ), .B0(n18136), .B1(
        \RAM<28><26> ), .Y(n2688) );
  AOI22X1 U1515 ( .A0(n18153), .A1(\RAM<27><26> ), .B0(n18150), .B1(
        \RAM<30><26> ), .Y(n2689) );
  AOI22X1 U1516 ( .A0(n18167), .A1(\RAM<29><26> ), .B0(n18164), .B1(
        \RAM<25><26> ), .Y(n2690) );
  NAND4X1 U1517 ( .A(n2634), .B(n2635), .C(n2636), .D(n2637), .Y(n2628) );
  AOI22X1 U1518 ( .A0(n18143), .A1(\RAM<47><27> ), .B0(n18136), .B1(
        \RAM<44><27> ), .Y(n2634) );
  AOI22X1 U1519 ( .A0(n18155), .A1(\RAM<43><27> ), .B0(n18150), .B1(
        \RAM<46><27> ), .Y(n2635) );
  AOI22X1 U1520 ( .A0(n2081), .A1(\RAM<45><27> ), .B0(n18164), .B1(
        \RAM<41><27> ), .Y(n2636) );
  NAND4X1 U1521 ( .A(n2624), .B(n2625), .C(n2626), .D(n2627), .Y(n2618) );
  AOI22X1 U1522 ( .A0(n18143), .A1(\RAM<63><27> ), .B0(n18136), .B1(
        \RAM<60><27> ), .Y(n2624) );
  AOI22X1 U1523 ( .A0(n18153), .A1(\RAM<59><27> ), .B0(n18150), .B1(
        \RAM<62><27> ), .Y(n2625) );
  AOI22X1 U1524 ( .A0(n18167), .A1(\RAM<61><27> ), .B0(n18164), .B1(
        \RAM<57><27> ), .Y(n2626) );
  NAND4X1 U1525 ( .A(n2644), .B(n2645), .C(n2646), .D(n2647), .Y(n2638) );
  AOI22X1 U1526 ( .A0(n18143), .A1(\RAM<31><27> ), .B0(n18136), .B1(
        \RAM<28><27> ), .Y(n2644) );
  AOI22X1 U1527 ( .A0(n18158), .A1(\RAM<27><27> ), .B0(n18150), .B1(
        \RAM<30><27> ), .Y(n2645) );
  AOI22X1 U1528 ( .A0(n18172), .A1(\RAM<29><27> ), .B0(n18164), .B1(
        \RAM<25><27> ), .Y(n2646) );
  NAND4X1 U1529 ( .A(n2580), .B(n2581), .C(n2582), .D(n2583), .Y(n2574) );
  AOI22X1 U1530 ( .A0(n18143), .A1(\RAM<63><28> ), .B0(n18136), .B1(
        \RAM<60><28> ), .Y(n2580) );
  AOI22X1 U1531 ( .A0(n18158), .A1(\RAM<59><28> ), .B0(n18150), .B1(
        \RAM<62><28> ), .Y(n2581) );
  AOI22X1 U1532 ( .A0(n18172), .A1(\RAM<61><28> ), .B0(n18164), .B1(
        \RAM<57><28> ), .Y(n2582) );
  NAND4X1 U1533 ( .A(n2590), .B(n2591), .C(n2592), .D(n2593), .Y(n2584) );
  AOI22X1 U1534 ( .A0(n18143), .A1(\RAM<47><28> ), .B0(n18136), .B1(
        \RAM<44><28> ), .Y(n2590) );
  AOI22X1 U1535 ( .A0(n18153), .A1(\RAM<43><28> ), .B0(n18150), .B1(
        \RAM<46><28> ), .Y(n2591) );
  AOI22X1 U1536 ( .A0(n18167), .A1(\RAM<45><28> ), .B0(n18164), .B1(
        \RAM<41><28> ), .Y(n2592) );
  NAND4X1 U1537 ( .A(n2600), .B(n2601), .C(n2602), .D(n2603), .Y(n2594) );
  AOI22X1 U1538 ( .A0(n18143), .A1(\RAM<31><28> ), .B0(n18136), .B1(
        \RAM<28><28> ), .Y(n2600) );
  AOI22X1 U1539 ( .A0(n18153), .A1(\RAM<27><28> ), .B0(n18150), .B1(
        \RAM<30><28> ), .Y(n2601) );
  AOI22X1 U1540 ( .A0(n18167), .A1(\RAM<29><28> ), .B0(n18164), .B1(
        \RAM<25><28> ), .Y(n2602) );
  NAND4X1 U1541 ( .A(n2536), .B(n2537), .C(n2538), .D(n2539), .Y(n2530) );
  AOI22X1 U1542 ( .A0(n18140), .A1(\RAM<63><29> ), .B0(n18137), .B1(
        \RAM<60><29> ), .Y(n2536) );
  AOI22X1 U1543 ( .A0(n18153), .A1(\RAM<59><29> ), .B0(n18151), .B1(
        \RAM<62><29> ), .Y(n2537) );
  AOI22X1 U1544 ( .A0(n18167), .A1(\RAM<61><29> ), .B0(n18165), .B1(
        \RAM<57><29> ), .Y(n2538) );
  NAND4X1 U1545 ( .A(n2546), .B(n2547), .C(n2548), .D(n2549), .Y(n2540) );
  AOI22X1 U1546 ( .A0(n18140), .A1(\RAM<47><29> ), .B0(n18134), .B1(
        \RAM<44><29> ), .Y(n2546) );
  AOI22X1 U1547 ( .A0(n18154), .A1(\RAM<43><29> ), .B0(n18148), .B1(
        \RAM<46><29> ), .Y(n2547) );
  AOI22X1 U1548 ( .A0(n18168), .A1(\RAM<45><29> ), .B0(n18162), .B1(
        \RAM<41><29> ), .Y(n2548) );
  NAND4X1 U1549 ( .A(n2556), .B(n2557), .C(n2558), .D(n2559), .Y(n2550) );
  AOI22X1 U1550 ( .A0(n18143), .A1(\RAM<31><29> ), .B0(n18134), .B1(
        \RAM<28><29> ), .Y(n2556) );
  AOI22X1 U1551 ( .A0(n2083), .A1(\RAM<27><29> ), .B0(n18148), .B1(
        \RAM<30><29> ), .Y(n2557) );
  AOI22X1 U1552 ( .A0(n2081), .A1(\RAM<29><29> ), .B0(n18162), .B1(
        \RAM<25><29> ), .Y(n2558) );
  NAND4X1 U1553 ( .A(n2458), .B(n2459), .C(n2460), .D(n2461), .Y(n2452) );
  AOI22X1 U1554 ( .A0(n18140), .A1(\RAM<47><30> ), .B0(n18137), .B1(
        \RAM<44><30> ), .Y(n2458) );
  AOI22X1 U1555 ( .A0(n18158), .A1(\RAM<43><30> ), .B0(n18149), .B1(
        \RAM<46><30> ), .Y(n2459) );
  AOI22X1 U1556 ( .A0(n18172), .A1(\RAM<45><30> ), .B0(n18163), .B1(
        \RAM<41><30> ), .Y(n2460) );
  NAND4X1 U1557 ( .A(n2448), .B(n2449), .C(n2450), .D(n2451), .Y(n2442) );
  AOI22X1 U1558 ( .A0(n18142), .A1(\RAM<63><30> ), .B0(n18135), .B1(
        \RAM<60><30> ), .Y(n2448) );
  AOI22X1 U1559 ( .A0(n18158), .A1(\RAM<59><30> ), .B0(n18149), .B1(
        \RAM<62><30> ), .Y(n2449) );
  AOI22X1 U1560 ( .A0(n18172), .A1(\RAM<61><30> ), .B0(n18163), .B1(
        \RAM<57><30> ), .Y(n2450) );
  NAND4X1 U1561 ( .A(n2468), .B(n2469), .C(n2470), .D(n2471), .Y(n2462) );
  AOI22X1 U1562 ( .A0(n18143), .A1(\RAM<31><30> ), .B0(n18134), .B1(
        \RAM<28><30> ), .Y(n2468) );
  AOI22X1 U1563 ( .A0(n2083), .A1(\RAM<27><30> ), .B0(n18148), .B1(
        \RAM<30><30> ), .Y(n2469) );
  AOI22X1 U1564 ( .A0(n2081), .A1(\RAM<29><30> ), .B0(n18162), .B1(
        \RAM<25><30> ), .Y(n2470) );
  NAND4X1 U1565 ( .A(n2394), .B(n2395), .C(n2396), .D(n2397), .Y(n2388) );
  AOI22X1 U1566 ( .A0(n2085), .A1(\RAM<15><31> ), .B0(n18132), .B1(
        \RAM<12><31> ), .Y(n2394) );
  AOI22X1 U1567 ( .A0(n18153), .A1(\RAM<11><31> ), .B0(n18146), .B1(
        \RAM<14><31> ), .Y(n2395) );
  AOI22X1 U1568 ( .A0(n18167), .A1(\RAM<13><31> ), .B0(n18164), .B1(
        \RAM<9><31> ), .Y(n2396) );
  NAND4X1 U1569 ( .A(n2404), .B(n2405), .C(n2406), .D(n2407), .Y(n2398) );
  AOI22X1 U1570 ( .A0(n18141), .A1(\RAM<63><31> ), .B0(n18133), .B1(
        \RAM<60><31> ), .Y(n2404) );
  AOI22X1 U1571 ( .A0(n18156), .A1(\RAM<59><31> ), .B0(n18150), .B1(
        \RAM<62><31> ), .Y(n2405) );
  AOI22X1 U1572 ( .A0(n18170), .A1(\RAM<61><31> ), .B0(n18164), .B1(
        \RAM<57><31> ), .Y(n2406) );
  NAND4X1 U1573 ( .A(n2424), .B(n2425), .C(n2426), .D(n2427), .Y(n2418) );
  AOI22X1 U1574 ( .A0(n18139), .A1(\RAM<31><31> ), .B0(n18132), .B1(
        \RAM<28><31> ), .Y(n2424) );
  AOI22X1 U1575 ( .A0(n18154), .A1(\RAM<27><31> ), .B0(n18147), .B1(
        \RAM<30><31> ), .Y(n2425) );
  AOI22X1 U1576 ( .A0(n18168), .A1(\RAM<29><31> ), .B0(n18161), .B1(
        \RAM<25><31> ), .Y(n2426) );
  NAND4X1 U1577 ( .A(n3450), .B(n3451), .C(n3452), .D(n3453), .Y(n3444) );
  AOI22X1 U1578 ( .A0(n18139), .A1(\RAM<15><0> ), .B0(n2086), .B1(\RAM<12><0> ), .Y(n3450) );
  AOI22X1 U1579 ( .A0(n18153), .A1(\RAM<11><0> ), .B0(n2084), .B1(\RAM<14><0> ), .Y(n3451) );
  AOI22X1 U1580 ( .A0(n18167), .A1(\RAM<13><0> ), .B0(n2082), .B1(\RAM<9><0> ), 
        .Y(n3452) );
  NAND4X1 U1581 ( .A(n3460), .B(n3461), .C(n3462), .D(n3463), .Y(n3454) );
  AOI22X1 U1582 ( .A0(n18139), .A1(\RAM<63><0> ), .B0(n18134), .B1(
        \RAM<60><0> ), .Y(n3460) );
  AOI22X1 U1583 ( .A0(n18153), .A1(\RAM<59><0> ), .B0(n18148), .B1(
        \RAM<62><0> ), .Y(n3461) );
  AOI22X1 U1584 ( .A0(n18167), .A1(\RAM<61><0> ), .B0(n18162), .B1(
        \RAM<57><0> ), .Y(n3462) );
  NAND4X1 U1585 ( .A(n3486), .B(n3487), .C(n3488), .D(n3489), .Y(n3474) );
  AOI22X1 U1586 ( .A0(n18139), .A1(\RAM<31><0> ), .B0(n18137), .B1(
        \RAM<28><0> ), .Y(n3486) );
  AOI22X1 U1587 ( .A0(n18153), .A1(\RAM<27><0> ), .B0(n18151), .B1(
        \RAM<30><0> ), .Y(n3487) );
  AOI22X1 U1588 ( .A0(n18167), .A1(\RAM<29><0> ), .B0(n18165), .B1(
        \RAM<25><0> ), .Y(n3488) );
  NAND4X1 U1589 ( .A(n2966), .B(n2967), .C(n2968), .D(n2969), .Y(n2960) );
  AOI22X1 U1590 ( .A0(n18143), .A1(\RAM<15><1> ), .B0(n18132), .B1(
        \RAM<12><1> ), .Y(n2966) );
  AOI22X1 U1591 ( .A0(n18156), .A1(\RAM<11><1> ), .B0(n18146), .B1(
        \RAM<14><1> ), .Y(n2967) );
  AOI22X1 U1592 ( .A0(n18170), .A1(\RAM<13><1> ), .B0(n18160), .B1(\RAM<9><1> ), .Y(n2968) );
  NAND4X1 U1593 ( .A(n2976), .B(n2977), .C(n2978), .D(n2979), .Y(n2970) );
  AOI22X1 U1594 ( .A0(n18140), .A1(\RAM<63><1> ), .B0(n18136), .B1(
        \RAM<60><1> ), .Y(n2976) );
  AOI22X1 U1595 ( .A0(n18156), .A1(\RAM<59><1> ), .B0(n18150), .B1(
        \RAM<62><1> ), .Y(n2977) );
  AOI22X1 U1596 ( .A0(n18170), .A1(\RAM<61><1> ), .B0(n18164), .B1(
        \RAM<57><1> ), .Y(n2978) );
  NAND4X1 U1597 ( .A(n2996), .B(n2997), .C(n2998), .D(n2999), .Y(n2990) );
  AOI22X1 U1598 ( .A0(n18143), .A1(\RAM<31><1> ), .B0(n18136), .B1(
        \RAM<28><1> ), .Y(n2996) );
  AOI22X1 U1599 ( .A0(n18156), .A1(\RAM<27><1> ), .B0(n18147), .B1(
        \RAM<30><1> ), .Y(n2997) );
  AOI22X1 U1600 ( .A0(n18170), .A1(\RAM<29><1> ), .B0(n18161), .B1(
        \RAM<25><1> ), .Y(n2998) );
  NAND4X1 U1601 ( .A(n2130), .B(n2131), .C(n2132), .D(n2133), .Y(n2124) );
  AOI22X1 U1602 ( .A0(n18139), .A1(\RAM<15><8> ), .B0(n18134), .B1(
        \RAM<12><8> ), .Y(n2130) );
  AOI22X1 U1603 ( .A0(n18153), .A1(\RAM<11><8> ), .B0(n18148), .B1(
        \RAM<14><8> ), .Y(n2131) );
  AOI22X1 U1604 ( .A0(n18167), .A1(\RAM<13><8> ), .B0(n18162), .B1(\RAM<9><8> ), .Y(n2132) );
  NAND4X1 U1605 ( .A(n2140), .B(n2141), .C(n2142), .D(n2143), .Y(n2134) );
  AOI22X1 U1606 ( .A0(n18141), .A1(\RAM<63><8> ), .B0(n18134), .B1(
        \RAM<60><8> ), .Y(n2140) );
  AOI22X1 U1607 ( .A0(n18155), .A1(\RAM<59><8> ), .B0(n18148), .B1(
        \RAM<62><8> ), .Y(n2141) );
  AOI22X1 U1608 ( .A0(n18169), .A1(\RAM<61><8> ), .B0(n18162), .B1(
        \RAM<57><8> ), .Y(n2142) );
  NAND4X1 U1609 ( .A(n2160), .B(n2161), .C(n2162), .D(n2163), .Y(n2154) );
  AOI22X1 U1610 ( .A0(n18141), .A1(\RAM<31><8> ), .B0(n18137), .B1(
        \RAM<28><8> ), .Y(n2160) );
  AOI22X1 U1611 ( .A0(n18157), .A1(\RAM<27><8> ), .B0(n18151), .B1(
        \RAM<30><8> ), .Y(n2161) );
  AOI22X1 U1612 ( .A0(n18171), .A1(\RAM<29><8> ), .B0(n18165), .B1(
        \RAM<25><8> ), .Y(n2162) );
  NAND4X1 U1613 ( .A(n2075), .B(n2076), .C(n2077), .D(n2078), .Y(n2060) );
  AOI22X1 U1614 ( .A0(n2085), .A1(\RAM<15><9> ), .B0(n18136), .B1(\RAM<12><9> ), .Y(n2075) );
  AOI22X1 U1615 ( .A0(n18154), .A1(\RAM<11><9> ), .B0(n18150), .B1(
        \RAM<14><9> ), .Y(n2076) );
  AOI22X1 U1616 ( .A0(n18168), .A1(\RAM<13><9> ), .B0(n18164), .B1(\RAM<9><9> ), .Y(n2077) );
  NAND4X1 U1617 ( .A(n2094), .B(n2095), .C(n2096), .D(n2097), .Y(n2087) );
  AOI22X1 U1618 ( .A0(n18144), .A1(\RAM<63><9> ), .B0(n18137), .B1(
        \RAM<60><9> ), .Y(n2094) );
  AOI22X1 U1619 ( .A0(n18158), .A1(\RAM<59><9> ), .B0(n18151), .B1(
        \RAM<62><9> ), .Y(n2095) );
  AOI22X1 U1620 ( .A0(n18172), .A1(\RAM<61><9> ), .B0(n18165), .B1(
        \RAM<57><9> ), .Y(n2096) );
  NAND4X1 U1621 ( .A(n2116), .B(n2117), .C(n2118), .D(n2119), .Y(n2109) );
  AOI22X1 U1622 ( .A0(n18144), .A1(\RAM<31><9> ), .B0(n18137), .B1(
        \RAM<28><9> ), .Y(n2116) );
  AOI22X1 U1623 ( .A0(n18157), .A1(\RAM<27><9> ), .B0(n18151), .B1(
        \RAM<30><9> ), .Y(n2117) );
  AOI22X1 U1624 ( .A0(n18171), .A1(\RAM<29><9> ), .B0(n18165), .B1(
        \RAM<25><9> ), .Y(n2118) );
  NAND4X1 U1625 ( .A(n2478), .B(n2479), .C(n2480), .D(n2481), .Y(n2477) );
  AOI22X1 U1626 ( .A0(n18199), .A1(\RAM<7><2> ), .B0(n18192), .B1(\RAM<4><2> ), 
        .Y(n2478) );
  AOI22X1 U1627 ( .A0(n2069), .A1(\RAM<5><2> ), .B0(n18220), .B1(\RAM<1><2> ), 
        .Y(n2480) );
  AOI22X1 U1628 ( .A0(n2071), .A1(\RAM<3><2> ), .B0(n18206), .B1(\RAM<6><2> ), 
        .Y(n2479) );
  NAND4X1 U1629 ( .A(n2488), .B(n2489), .C(n2490), .D(n2491), .Y(n2487) );
  AOI22X1 U1630 ( .A0(n18199), .A1(\RAM<55><2> ), .B0(n2074), .B1(\RAM<52><2> ), .Y(n2488) );
  AOI22X1 U1631 ( .A0(n2069), .A1(\RAM<53><2> ), .B0(n18220), .B1(\RAM<49><2> ), .Y(n2490) );
  AOI22X1 U1632 ( .A0(n18209), .A1(\RAM<51><2> ), .B0(n18206), .B1(
        \RAM<54><2> ), .Y(n2489) );
  NAND4X1 U1633 ( .A(n2508), .B(n2509), .C(n2510), .D(n2511), .Y(n2507) );
  AOI22X1 U1634 ( .A0(n18197), .A1(\RAM<23><2> ), .B0(n2074), .B1(\RAM<20><2> ), .Y(n2508) );
  AOI22X1 U1635 ( .A0(n18227), .A1(\RAM<21><2> ), .B0(n18220), .B1(
        \RAM<17><2> ), .Y(n2510) );
  AOI22X1 U1636 ( .A0(n18209), .A1(\RAM<19><2> ), .B0(n18206), .B1(
        \RAM<22><2> ), .Y(n2509) );
  NAND4X1 U1637 ( .A(n2346), .B(n2347), .C(n2348), .D(n2349), .Y(n2345) );
  AOI22X1 U1638 ( .A0(n18196), .A1(\RAM<7><3> ), .B0(n18192), .B1(\RAM<4><3> ), 
        .Y(n2346) );
  AOI22X1 U1639 ( .A0(n18225), .A1(\RAM<5><3> ), .B0(n18220), .B1(\RAM<1><3> ), 
        .Y(n2348) );
  AOI22X1 U1640 ( .A0(n18212), .A1(\RAM<3><3> ), .B0(n18203), .B1(\RAM<6><3> ), 
        .Y(n2347) );
  NAND4X1 U1641 ( .A(n2356), .B(n2357), .C(n2358), .D(n2359), .Y(n2355) );
  AOI22X1 U1642 ( .A0(n18195), .A1(\RAM<55><3> ), .B0(n18192), .B1(
        \RAM<52><3> ), .Y(n2356) );
  AOI22X1 U1643 ( .A0(n18225), .A1(\RAM<53><3> ), .B0(n18218), .B1(
        \RAM<49><3> ), .Y(n2358) );
  AOI22X1 U1644 ( .A0(n18212), .A1(\RAM<51><3> ), .B0(n18204), .B1(
        \RAM<54><3> ), .Y(n2357) );
  NAND4X1 U1645 ( .A(n2376), .B(n2377), .C(n2378), .D(n2379), .Y(n2375) );
  AOI22X1 U1646 ( .A0(n18200), .A1(\RAM<23><3> ), .B0(n18192), .B1(
        \RAM<20><3> ), .Y(n2376) );
  AOI22X1 U1647 ( .A0(n18224), .A1(\RAM<21><3> ), .B0(n18218), .B1(
        \RAM<17><3> ), .Y(n2378) );
  AOI22X1 U1648 ( .A0(n18212), .A1(\RAM<19><3> ), .B0(n18203), .B1(
        \RAM<22><3> ), .Y(n2377) );
  NAND4X1 U1649 ( .A(n2302), .B(n2303), .C(n2304), .D(n2305), .Y(n2301) );
  AOI22X1 U1650 ( .A0(n18195), .A1(\RAM<7><4> ), .B0(n18192), .B1(\RAM<4><4> ), 
        .Y(n2302) );
  AOI22X1 U1651 ( .A0(n18228), .A1(\RAM<5><4> ), .B0(n18218), .B1(\RAM<1><4> ), 
        .Y(n2304) );
  AOI22X1 U1652 ( .A0(n2071), .A1(\RAM<3><4> ), .B0(n18204), .B1(\RAM<6><4> ), 
        .Y(n2303) );
  NAND4X1 U1653 ( .A(n2312), .B(n2313), .C(n2314), .D(n2315), .Y(n2311) );
  AOI22X1 U1654 ( .A0(n18196), .A1(\RAM<55><4> ), .B0(n18192), .B1(
        \RAM<52><4> ), .Y(n2312) );
  AOI22X1 U1655 ( .A0(n18224), .A1(\RAM<53><4> ), .B0(n18220), .B1(
        \RAM<49><4> ), .Y(n2314) );
  AOI22X1 U1656 ( .A0(n18212), .A1(\RAM<51><4> ), .B0(n18203), .B1(
        \RAM<54><4> ), .Y(n2313) );
  NAND4X1 U1657 ( .A(n2332), .B(n2333), .C(n2334), .D(n2335), .Y(n2331) );
  AOI22X1 U1658 ( .A0(n18196), .A1(\RAM<23><4> ), .B0(n18192), .B1(
        \RAM<20><4> ), .Y(n2332) );
  AOI22X1 U1659 ( .A0(n18224), .A1(\RAM<21><4> ), .B0(n18220), .B1(
        \RAM<17><4> ), .Y(n2334) );
  AOI22X1 U1660 ( .A0(n18213), .A1(\RAM<19><4> ), .B0(n18202), .B1(
        \RAM<22><4> ), .Y(n2333) );
  NAND4X1 U1661 ( .A(n2258), .B(n2259), .C(n2260), .D(n2261), .Y(n2257) );
  AOI22X1 U1662 ( .A0(n18200), .A1(\RAM<7><5> ), .B0(n18193), .B1(\RAM<4><5> ), 
        .Y(n2258) );
  AOI22X1 U1663 ( .A0(n18228), .A1(\RAM<5><5> ), .B0(n18221), .B1(\RAM<1><5> ), 
        .Y(n2260) );
  AOI22X1 U1664 ( .A0(n2071), .A1(\RAM<3><5> ), .B0(n18207), .B1(\RAM<6><5> ), 
        .Y(n2259) );
  NAND4X1 U1665 ( .A(n2268), .B(n2269), .C(n2270), .D(n2271), .Y(n2267) );
  AOI22X1 U1666 ( .A0(n18200), .A1(\RAM<55><5> ), .B0(n18193), .B1(
        \RAM<52><5> ), .Y(n2268) );
  AOI22X1 U1667 ( .A0(n18228), .A1(\RAM<53><5> ), .B0(n18221), .B1(
        \RAM<49><5> ), .Y(n2270) );
  AOI22X1 U1668 ( .A0(n18214), .A1(\RAM<51><5> ), .B0(n18207), .B1(
        \RAM<54><5> ), .Y(n2269) );
  NAND4X1 U1669 ( .A(n2288), .B(n2289), .C(n2290), .D(n2291), .Y(n2287) );
  AOI22X1 U1670 ( .A0(n18200), .A1(\RAM<23><5> ), .B0(n18193), .B1(
        \RAM<20><5> ), .Y(n2288) );
  AOI22X1 U1671 ( .A0(n18228), .A1(\RAM<21><5> ), .B0(n18221), .B1(
        \RAM<17><5> ), .Y(n2290) );
  AOI22X1 U1672 ( .A0(n18211), .A1(\RAM<19><5> ), .B0(n18207), .B1(
        \RAM<22><5> ), .Y(n2289) );
  NAND4X1 U1673 ( .A(n2214), .B(n2215), .C(n2216), .D(n2217), .Y(n2213) );
  AOI22X1 U1674 ( .A0(n18200), .A1(\RAM<7><6> ), .B0(n18193), .B1(\RAM<4><6> ), 
        .Y(n2214) );
  AOI22X1 U1675 ( .A0(n18228), .A1(\RAM<5><6> ), .B0(n18221), .B1(\RAM<1><6> ), 
        .Y(n2216) );
  AOI22X1 U1676 ( .A0(n2071), .A1(\RAM<3><6> ), .B0(n18207), .B1(\RAM<6><6> ), 
        .Y(n2215) );
  NAND4X1 U1677 ( .A(n2224), .B(n2225), .C(n2226), .D(n2227), .Y(n2223) );
  AOI22X1 U1678 ( .A0(n18200), .A1(\RAM<55><6> ), .B0(n18193), .B1(
        \RAM<52><6> ), .Y(n2224) );
  AOI22X1 U1679 ( .A0(n18228), .A1(\RAM<53><6> ), .B0(n18221), .B1(
        \RAM<49><6> ), .Y(n2226) );
  AOI22X1 U1680 ( .A0(n18211), .A1(\RAM<51><6> ), .B0(n18207), .B1(
        \RAM<54><6> ), .Y(n2225) );
  NAND4X1 U1681 ( .A(n2244), .B(n2245), .C(n2246), .D(n2247), .Y(n2243) );
  AOI22X1 U1682 ( .A0(n18200), .A1(\RAM<23><6> ), .B0(n18193), .B1(
        \RAM<20><6> ), .Y(n2244) );
  AOI22X1 U1683 ( .A0(n18228), .A1(\RAM<21><6> ), .B0(n18221), .B1(
        \RAM<17><6> ), .Y(n2246) );
  AOI22X1 U1684 ( .A0(n18210), .A1(\RAM<19><6> ), .B0(n18207), .B1(
        \RAM<22><6> ), .Y(n2245) );
  NAND4X1 U1685 ( .A(n2170), .B(n2171), .C(n2172), .D(n2173), .Y(n2169) );
  AOI22X1 U1686 ( .A0(n18200), .A1(\RAM<7><7> ), .B0(n18193), .B1(\RAM<4><7> ), 
        .Y(n2170) );
  AOI22X1 U1687 ( .A0(n18228), .A1(\RAM<5><7> ), .B0(n18221), .B1(\RAM<1><7> ), 
        .Y(n2172) );
  AOI22X1 U1688 ( .A0(n2071), .A1(\RAM<3><7> ), .B0(n18207), .B1(\RAM<6><7> ), 
        .Y(n2171) );
  NAND4X1 U1689 ( .A(n2180), .B(n2181), .C(n2182), .D(n2183), .Y(n2179) );
  AOI22X1 U1690 ( .A0(n18200), .A1(\RAM<55><7> ), .B0(n18193), .B1(
        \RAM<52><7> ), .Y(n2180) );
  AOI22X1 U1691 ( .A0(n18228), .A1(\RAM<53><7> ), .B0(n18221), .B1(
        \RAM<49><7> ), .Y(n2182) );
  AOI22X1 U1692 ( .A0(n18210), .A1(\RAM<51><7> ), .B0(n18207), .B1(
        \RAM<54><7> ), .Y(n2181) );
  NAND4X1 U1693 ( .A(n2200), .B(n2201), .C(n2202), .D(n2203), .Y(n2199) );
  AOI22X1 U1694 ( .A0(n18200), .A1(\RAM<23><7> ), .B0(n18193), .B1(
        \RAM<20><7> ), .Y(n2200) );
  AOI22X1 U1695 ( .A0(n18228), .A1(\RAM<21><7> ), .B0(n18221), .B1(
        \RAM<17><7> ), .Y(n2202) );
  AOI22X1 U1696 ( .A0(n18214), .A1(\RAM<19><7> ), .B0(n18207), .B1(
        \RAM<22><7> ), .Y(n2201) );
  NAND4X1 U1697 ( .A(n3402), .B(n3403), .C(n3404), .D(n3405), .Y(n3401) );
  AOI22X1 U1698 ( .A0(n2073), .A1(\RAM<7><10> ), .B0(n18188), .B1(\RAM<4><10> ), .Y(n3402) );
  AOI22X1 U1699 ( .A0(n18227), .A1(\RAM<5><10> ), .B0(n18220), .B1(
        \RAM<1><10> ), .Y(n3404) );
  AOI22X1 U1700 ( .A0(n18209), .A1(\RAM<3><10> ), .B0(n18206), .B1(
        \RAM<6><10> ), .Y(n3403) );
  NAND4X1 U1701 ( .A(n3412), .B(n3413), .C(n3414), .D(n3415), .Y(n3411) );
  AOI22X1 U1702 ( .A0(n18197), .A1(\RAM<55><10> ), .B0(n18188), .B1(
        \RAM<52><10> ), .Y(n3412) );
  AOI22X1 U1703 ( .A0(n18228), .A1(\RAM<53><10> ), .B0(n18219), .B1(
        \RAM<49><10> ), .Y(n3414) );
  AOI22X1 U1704 ( .A0(n18209), .A1(\RAM<51><10> ), .B0(n18207), .B1(
        \RAM<54><10> ), .Y(n3413) );
  NAND4X1 U1705 ( .A(n3432), .B(n3433), .C(n3434), .D(n3435), .Y(n3431) );
  AOI22X1 U1706 ( .A0(n18199), .A1(\RAM<23><10> ), .B0(n18188), .B1(
        \RAM<20><10> ), .Y(n3432) );
  AOI22X1 U1707 ( .A0(n18228), .A1(\RAM<21><10> ), .B0(n18218), .B1(
        \RAM<17><10> ), .Y(n3434) );
  AOI22X1 U1708 ( .A0(n18209), .A1(\RAM<19><10> ), .B0(n18207), .B1(
        \RAM<22><10> ), .Y(n3433) );
  NAND4X1 U1709 ( .A(n3358), .B(n3359), .C(n3360), .D(n3361), .Y(n3357) );
  AOI22X1 U1710 ( .A0(n18196), .A1(\RAM<7><11> ), .B0(n18188), .B1(
        \RAM<4><11> ), .Y(n3358) );
  AOI22X1 U1711 ( .A0(n18225), .A1(\RAM<5><11> ), .B0(n18219), .B1(
        \RAM<1><11> ), .Y(n3360) );
  AOI22X1 U1712 ( .A0(n18209), .A1(\RAM<3><11> ), .B0(n18205), .B1(
        \RAM<6><11> ), .Y(n3359) );
  NAND4X1 U1713 ( .A(n3368), .B(n3369), .C(n3370), .D(n3371), .Y(n3367) );
  AOI22X1 U1714 ( .A0(n18199), .A1(\RAM<55><11> ), .B0(n18188), .B1(
        \RAM<52><11> ), .Y(n3368) );
  AOI22X1 U1715 ( .A0(n18228), .A1(\RAM<53><11> ), .B0(n18218), .B1(
        \RAM<49><11> ), .Y(n3370) );
  AOI22X1 U1716 ( .A0(n18209), .A1(\RAM<51><11> ), .B0(n18206), .B1(
        \RAM<54><11> ), .Y(n3369) );
  NAND4X1 U1717 ( .A(n3388), .B(n3389), .C(n3390), .D(n3391), .Y(n3387) );
  AOI22X1 U1718 ( .A0(n18198), .A1(\RAM<23><11> ), .B0(n18188), .B1(
        \RAM<20><11> ), .Y(n3388) );
  AOI22X1 U1719 ( .A0(n18226), .A1(\RAM<21><11> ), .B0(n18220), .B1(
        \RAM<17><11> ), .Y(n3390) );
  AOI22X1 U1720 ( .A0(n18209), .A1(\RAM<19><11> ), .B0(n18206), .B1(
        \RAM<22><11> ), .Y(n3389) );
  NAND4X1 U1721 ( .A(n3334), .B(n3335), .C(n3336), .D(n3337), .Y(n3333) );
  AOI22X1 U1722 ( .A0(n18195), .A1(\RAM<39><12> ), .B0(n18189), .B1(
        \RAM<36><12> ), .Y(n3334) );
  AOI22X1 U1723 ( .A0(n18223), .A1(\RAM<37><12> ), .B0(n18216), .B1(
        \RAM<33><12> ), .Y(n3336) );
  AOI22X1 U1724 ( .A0(n18210), .A1(\RAM<35><12> ), .B0(n18202), .B1(
        \RAM<38><12> ), .Y(n3335) );
  NAND4X1 U1725 ( .A(n3324), .B(n3325), .C(n3326), .D(n3327), .Y(n3323) );
  AOI22X1 U1726 ( .A0(n18195), .A1(\RAM<55><12> ), .B0(n18189), .B1(
        \RAM<52><12> ), .Y(n3324) );
  AOI22X1 U1727 ( .A0(n18223), .A1(\RAM<53><12> ), .B0(n18216), .B1(
        \RAM<49><12> ), .Y(n3326) );
  AOI22X1 U1728 ( .A0(n18210), .A1(\RAM<51><12> ), .B0(n18202), .B1(
        \RAM<54><12> ), .Y(n3325) );
  NAND4X1 U1729 ( .A(n3344), .B(n3345), .C(n3346), .D(n3347), .Y(n3343) );
  AOI22X1 U1730 ( .A0(n18195), .A1(\RAM<23><12> ), .B0(n18189), .B1(
        \RAM<20><12> ), .Y(n3344) );
  AOI22X1 U1731 ( .A0(n18223), .A1(\RAM<21><12> ), .B0(n18216), .B1(
        \RAM<17><12> ), .Y(n3346) );
  AOI22X1 U1732 ( .A0(n18210), .A1(\RAM<19><12> ), .B0(n18202), .B1(
        \RAM<22><12> ), .Y(n3345) );
  NAND4X1 U1733 ( .A(n3290), .B(n3291), .C(n3292), .D(n3293), .Y(n3289) );
  AOI22X1 U1734 ( .A0(n18195), .A1(\RAM<39><13> ), .B0(n18189), .B1(
        \RAM<36><13> ), .Y(n3290) );
  AOI22X1 U1735 ( .A0(n18223), .A1(\RAM<37><13> ), .B0(n18216), .B1(
        \RAM<33><13> ), .Y(n3292) );
  AOI22X1 U1736 ( .A0(n18210), .A1(\RAM<35><13> ), .B0(n18202), .B1(
        \RAM<38><13> ), .Y(n3291) );
  NAND4X1 U1737 ( .A(n3280), .B(n3281), .C(n3282), .D(n3283), .Y(n3279) );
  AOI22X1 U1738 ( .A0(n18195), .A1(\RAM<55><13> ), .B0(n18189), .B1(
        \RAM<52><13> ), .Y(n3280) );
  AOI22X1 U1739 ( .A0(n18223), .A1(\RAM<53><13> ), .B0(n18216), .B1(
        \RAM<49><13> ), .Y(n3282) );
  AOI22X1 U1740 ( .A0(n18210), .A1(\RAM<51><13> ), .B0(n18202), .B1(
        \RAM<54><13> ), .Y(n3281) );
  NAND4X1 U1741 ( .A(n3300), .B(n3301), .C(n3302), .D(n3303), .Y(n3299) );
  AOI22X1 U1742 ( .A0(n18195), .A1(\RAM<23><13> ), .B0(n18189), .B1(
        \RAM<20><13> ), .Y(n3300) );
  AOI22X1 U1743 ( .A0(n18223), .A1(\RAM<21><13> ), .B0(n18216), .B1(
        \RAM<17><13> ), .Y(n3302) );
  AOI22X1 U1744 ( .A0(n18210), .A1(\RAM<19><13> ), .B0(n18202), .B1(
        \RAM<22><13> ), .Y(n3301) );
  NAND4X1 U1745 ( .A(n3246), .B(n3247), .C(n3248), .D(n3249), .Y(n3245) );
  AOI22X1 U1746 ( .A0(n18195), .A1(\RAM<39><14> ), .B0(n18189), .B1(
        \RAM<36><14> ), .Y(n3246) );
  AOI22X1 U1747 ( .A0(n18223), .A1(\RAM<37><14> ), .B0(n18216), .B1(
        \RAM<33><14> ), .Y(n3248) );
  AOI22X1 U1748 ( .A0(n18210), .A1(\RAM<35><14> ), .B0(n18202), .B1(
        \RAM<38><14> ), .Y(n3247) );
  NAND4X1 U1749 ( .A(n3236), .B(n3237), .C(n3238), .D(n3239), .Y(n3235) );
  AOI22X1 U1750 ( .A0(n18195), .A1(\RAM<55><14> ), .B0(n18189), .B1(
        \RAM<52><14> ), .Y(n3236) );
  AOI22X1 U1751 ( .A0(n18223), .A1(\RAM<53><14> ), .B0(n18216), .B1(
        \RAM<49><14> ), .Y(n3238) );
  AOI22X1 U1752 ( .A0(n18210), .A1(\RAM<51><14> ), .B0(n18202), .B1(
        \RAM<54><14> ), .Y(n3237) );
  NAND4X1 U1753 ( .A(n3256), .B(n3257), .C(n3258), .D(n3259), .Y(n3255) );
  AOI22X1 U1754 ( .A0(n18195), .A1(\RAM<23><14> ), .B0(n18189), .B1(
        \RAM<20><14> ), .Y(n3256) );
  AOI22X1 U1755 ( .A0(n18223), .A1(\RAM<21><14> ), .B0(n18216), .B1(
        \RAM<17><14> ), .Y(n3258) );
  AOI22X1 U1756 ( .A0(n18210), .A1(\RAM<19><14> ), .B0(n18202), .B1(
        \RAM<22><14> ), .Y(n3257) );
  NAND4X1 U1757 ( .A(n3202), .B(n3203), .C(n3204), .D(n3205), .Y(n3201) );
  AOI22X1 U1758 ( .A0(n18196), .A1(\RAM<39><15> ), .B0(n18190), .B1(
        \RAM<36><15> ), .Y(n3202) );
  AOI22X1 U1759 ( .A0(n18224), .A1(\RAM<37><15> ), .B0(n18217), .B1(
        \RAM<33><15> ), .Y(n3204) );
  AOI22X1 U1760 ( .A0(n18211), .A1(\RAM<35><15> ), .B0(n18203), .B1(
        \RAM<38><15> ), .Y(n3203) );
  NAND4X1 U1761 ( .A(n3192), .B(n3193), .C(n3194), .D(n3195), .Y(n3191) );
  AOI22X1 U1762 ( .A0(n18196), .A1(\RAM<55><15> ), .B0(n18190), .B1(
        \RAM<52><15> ), .Y(n3192) );
  AOI22X1 U1763 ( .A0(n18224), .A1(\RAM<53><15> ), .B0(n18217), .B1(
        \RAM<49><15> ), .Y(n3194) );
  AOI22X1 U1764 ( .A0(n18211), .A1(\RAM<51><15> ), .B0(n18203), .B1(
        \RAM<54><15> ), .Y(n3193) );
  NAND4X1 U1765 ( .A(n3212), .B(n3213), .C(n3214), .D(n3215), .Y(n3211) );
  AOI22X1 U1766 ( .A0(n18196), .A1(\RAM<23><15> ), .B0(n18190), .B1(
        \RAM<20><15> ), .Y(n3212) );
  AOI22X1 U1767 ( .A0(n18224), .A1(\RAM<21><15> ), .B0(n18217), .B1(
        \RAM<17><15> ), .Y(n3214) );
  AOI22X1 U1768 ( .A0(n18211), .A1(\RAM<19><15> ), .B0(n18203), .B1(
        \RAM<22><15> ), .Y(n3213) );
  NAND4X1 U1769 ( .A(n3138), .B(n3139), .C(n3140), .D(n3141), .Y(n3137) );
  AOI22X1 U1770 ( .A0(n18196), .A1(\RAM<7><16> ), .B0(n18190), .B1(
        \RAM<4><16> ), .Y(n3138) );
  AOI22X1 U1771 ( .A0(n18224), .A1(\RAM<5><16> ), .B0(n18217), .B1(
        \RAM<1><16> ), .Y(n3140) );
  AOI22X1 U1772 ( .A0(n18211), .A1(\RAM<3><16> ), .B0(n18203), .B1(
        \RAM<6><16> ), .Y(n3139) );
  NAND4X1 U1773 ( .A(n3148), .B(n3149), .C(n3150), .D(n3151), .Y(n3147) );
  AOI22X1 U1774 ( .A0(n18196), .A1(\RAM<55><16> ), .B0(n18190), .B1(
        \RAM<52><16> ), .Y(n3148) );
  AOI22X1 U1775 ( .A0(n18224), .A1(\RAM<53><16> ), .B0(n18217), .B1(
        \RAM<49><16> ), .Y(n3150) );
  AOI22X1 U1776 ( .A0(n18211), .A1(\RAM<51><16> ), .B0(n18203), .B1(
        \RAM<54><16> ), .Y(n3149) );
  NAND4X1 U1777 ( .A(n3168), .B(n3169), .C(n3170), .D(n3171), .Y(n3167) );
  AOI22X1 U1778 ( .A0(n18196), .A1(\RAM<23><16> ), .B0(n18190), .B1(
        \RAM<20><16> ), .Y(n3168) );
  AOI22X1 U1779 ( .A0(n18224), .A1(\RAM<21><16> ), .B0(n18217), .B1(
        \RAM<17><16> ), .Y(n3170) );
  AOI22X1 U1780 ( .A0(n18211), .A1(\RAM<19><16> ), .B0(n18203), .B1(
        \RAM<22><16> ), .Y(n3169) );
  NAND4X1 U1781 ( .A(n3094), .B(n3095), .C(n3096), .D(n3097), .Y(n3093) );
  AOI22X1 U1782 ( .A0(n18196), .A1(\RAM<7><17> ), .B0(n18190), .B1(
        \RAM<4><17> ), .Y(n3094) );
  AOI22X1 U1783 ( .A0(n18224), .A1(\RAM<5><17> ), .B0(n18217), .B1(
        \RAM<1><17> ), .Y(n3096) );
  AOI22X1 U1784 ( .A0(n18211), .A1(\RAM<3><17> ), .B0(n18203), .B1(
        \RAM<6><17> ), .Y(n3095) );
  NAND4X1 U1785 ( .A(n3104), .B(n3105), .C(n3106), .D(n3107), .Y(n3103) );
  AOI22X1 U1786 ( .A0(n18196), .A1(\RAM<55><17> ), .B0(n18190), .B1(
        \RAM<52><17> ), .Y(n3104) );
  AOI22X1 U1787 ( .A0(n18224), .A1(\RAM<53><17> ), .B0(n18217), .B1(
        \RAM<49><17> ), .Y(n3106) );
  AOI22X1 U1788 ( .A0(n18211), .A1(\RAM<51><17> ), .B0(n18203), .B1(
        \RAM<54><17> ), .Y(n3105) );
  NAND4X1 U1789 ( .A(n3124), .B(n3125), .C(n3126), .D(n3127), .Y(n3123) );
  AOI22X1 U1790 ( .A0(n18196), .A1(\RAM<23><17> ), .B0(n18190), .B1(
        \RAM<20><17> ), .Y(n3124) );
  AOI22X1 U1791 ( .A0(n18224), .A1(\RAM<21><17> ), .B0(n18217), .B1(
        \RAM<17><17> ), .Y(n3126) );
  AOI22X1 U1792 ( .A0(n18211), .A1(\RAM<19><17> ), .B0(n18203), .B1(
        \RAM<22><17> ), .Y(n3125) );
  NAND4X1 U1793 ( .A(n3050), .B(n3051), .C(n3052), .D(n3053), .Y(n3049) );
  AOI22X1 U1794 ( .A0(n2073), .A1(\RAM<7><18> ), .B0(n18189), .B1(\RAM<4><18> ), .Y(n3050) );
  AOI22X1 U1795 ( .A0(n2069), .A1(\RAM<5><18> ), .B0(n18217), .B1(\RAM<1><18> ), .Y(n3052) );
  AOI22X1 U1796 ( .A0(n18211), .A1(\RAM<3><18> ), .B0(n18204), .B1(
        \RAM<6><18> ), .Y(n3051) );
  NAND4X1 U1797 ( .A(n3060), .B(n3061), .C(n3062), .D(n3063), .Y(n3059) );
  AOI22X1 U1798 ( .A0(n2073), .A1(\RAM<55><18> ), .B0(n18193), .B1(
        \RAM<52><18> ), .Y(n3060) );
  AOI22X1 U1799 ( .A0(n18224), .A1(\RAM<53><18> ), .B0(n18217), .B1(
        \RAM<49><18> ), .Y(n3062) );
  AOI22X1 U1800 ( .A0(n18211), .A1(\RAM<51><18> ), .B0(n18204), .B1(
        \RAM<54><18> ), .Y(n3061) );
  NAND4X1 U1801 ( .A(n3080), .B(n3081), .C(n3082), .D(n3083), .Y(n3079) );
  AOI22X1 U1802 ( .A0(n18195), .A1(\RAM<23><18> ), .B0(n18190), .B1(
        \RAM<20><18> ), .Y(n3080) );
  AOI22X1 U1803 ( .A0(n18223), .A1(\RAM<21><18> ), .B0(n18217), .B1(
        \RAM<17><18> ), .Y(n3082) );
  AOI22X1 U1804 ( .A0(n18211), .A1(\RAM<19><18> ), .B0(n18203), .B1(
        \RAM<22><18> ), .Y(n3081) );
  NAND4X1 U1805 ( .A(n3006), .B(n3007), .C(n3008), .D(n3009), .Y(n3005) );
  AOI22X1 U1806 ( .A0(n2073), .A1(\RAM<7><19> ), .B0(n18188), .B1(\RAM<4><19> ), .Y(n3006) );
  AOI22X1 U1807 ( .A0(n2069), .A1(\RAM<5><19> ), .B0(n18216), .B1(\RAM<1><19> ), .Y(n3008) );
  AOI22X1 U1808 ( .A0(n18210), .A1(\RAM<3><19> ), .B0(n2072), .B1(\RAM<6><19> ), .Y(n3007) );
  NAND4X1 U1809 ( .A(n3016), .B(n3017), .C(n3018), .D(n3019), .Y(n3015) );
  AOI22X1 U1810 ( .A0(n2073), .A1(\RAM<55><19> ), .B0(n18190), .B1(
        \RAM<52><19> ), .Y(n3016) );
  AOI22X1 U1811 ( .A0(n18223), .A1(\RAM<53><19> ), .B0(n18216), .B1(
        \RAM<49><19> ), .Y(n3018) );
  AOI22X1 U1812 ( .A0(n18210), .A1(\RAM<51><19> ), .B0(n18203), .B1(
        \RAM<54><19> ), .Y(n3017) );
  NAND4X1 U1813 ( .A(n3036), .B(n3037), .C(n3038), .D(n3039), .Y(n3035) );
  AOI22X1 U1814 ( .A0(n18200), .A1(\RAM<23><19> ), .B0(n18189), .B1(
        \RAM<20><19> ), .Y(n3036) );
  AOI22X1 U1815 ( .A0(n18225), .A1(\RAM<21><19> ), .B0(n18216), .B1(
        \RAM<17><19> ), .Y(n3038) );
  AOI22X1 U1816 ( .A0(n18210), .A1(\RAM<19><19> ), .B0(n18202), .B1(
        \RAM<22><19> ), .Y(n3037) );
  NAND4X1 U1817 ( .A(n2938), .B(n2939), .C(n2940), .D(n2941), .Y(n2937) );
  AOI22X1 U1818 ( .A0(n18197), .A1(\RAM<39><20> ), .B0(n2074), .B1(
        \RAM<36><20> ), .Y(n2938) );
  AOI22X1 U1819 ( .A0(n18225), .A1(\RAM<37><20> ), .B0(n18218), .B1(
        \RAM<33><20> ), .Y(n2940) );
  AOI22X1 U1820 ( .A0(n18212), .A1(\RAM<35><20> ), .B0(n18204), .B1(
        \RAM<38><20> ), .Y(n2939) );
  NAND4X1 U1821 ( .A(n2928), .B(n2929), .C(n2930), .D(n2931), .Y(n2927) );
  AOI22X1 U1822 ( .A0(n18197), .A1(\RAM<55><20> ), .B0(n2074), .B1(
        \RAM<52><20> ), .Y(n2928) );
  AOI22X1 U1823 ( .A0(n18225), .A1(\RAM<53><20> ), .B0(n18218), .B1(
        \RAM<49><20> ), .Y(n2930) );
  AOI22X1 U1824 ( .A0(n18212), .A1(\RAM<51><20> ), .B0(n18204), .B1(
        \RAM<54><20> ), .Y(n2929) );
  NAND4X1 U1825 ( .A(n2948), .B(n2949), .C(n2950), .D(n2951), .Y(n2947) );
  AOI22X1 U1826 ( .A0(n18197), .A1(\RAM<23><20> ), .B0(n18189), .B1(
        \RAM<20><20> ), .Y(n2948) );
  AOI22X1 U1827 ( .A0(n18225), .A1(\RAM<21><20> ), .B0(n18218), .B1(
        \RAM<17><20> ), .Y(n2950) );
  AOI22X1 U1828 ( .A0(n18212), .A1(\RAM<19><20> ), .B0(n18204), .B1(
        \RAM<22><20> ), .Y(n2949) );
  NAND4X1 U1829 ( .A(n2874), .B(n2875), .C(n2876), .D(n2877), .Y(n2873) );
  AOI22X1 U1830 ( .A0(n18197), .A1(\RAM<7><21> ), .B0(n18193), .B1(
        \RAM<4><21> ), .Y(n2874) );
  AOI22X1 U1831 ( .A0(n18225), .A1(\RAM<5><21> ), .B0(n18218), .B1(
        \RAM<1><21> ), .Y(n2876) );
  AOI22X1 U1832 ( .A0(n18212), .A1(\RAM<3><21> ), .B0(n18204), .B1(
        \RAM<6><21> ), .Y(n2875) );
  NAND4X1 U1833 ( .A(n2884), .B(n2885), .C(n2886), .D(n2887), .Y(n2883) );
  AOI22X1 U1834 ( .A0(n18197), .A1(\RAM<55><21> ), .B0(n2074), .B1(
        \RAM<52><21> ), .Y(n2884) );
  AOI22X1 U1835 ( .A0(n18225), .A1(\RAM<53><21> ), .B0(n18218), .B1(
        \RAM<49><21> ), .Y(n2886) );
  AOI22X1 U1836 ( .A0(n18212), .A1(\RAM<51><21> ), .B0(n18204), .B1(
        \RAM<54><21> ), .Y(n2885) );
  NAND4X1 U1837 ( .A(n2904), .B(n2905), .C(n2906), .D(n2907), .Y(n2903) );
  AOI22X1 U1838 ( .A0(n18197), .A1(\RAM<23><21> ), .B0(n18189), .B1(
        \RAM<20><21> ), .Y(n2904) );
  AOI22X1 U1839 ( .A0(n18225), .A1(\RAM<21><21> ), .B0(n18218), .B1(
        \RAM<17><21> ), .Y(n2906) );
  AOI22X1 U1840 ( .A0(n18212), .A1(\RAM<19><21> ), .B0(n18204), .B1(
        \RAM<22><21> ), .Y(n2905) );
  NAND4X1 U1841 ( .A(n2830), .B(n2831), .C(n2832), .D(n2833), .Y(n2829) );
  AOI22X1 U1842 ( .A0(n18197), .A1(\RAM<7><22> ), .B0(n18190), .B1(
        \RAM<4><22> ), .Y(n2830) );
  AOI22X1 U1843 ( .A0(n18225), .A1(\RAM<5><22> ), .B0(n18218), .B1(
        \RAM<1><22> ), .Y(n2832) );
  AOI22X1 U1844 ( .A0(n18212), .A1(\RAM<3><22> ), .B0(n18204), .B1(
        \RAM<6><22> ), .Y(n2831) );
  NAND4X1 U1845 ( .A(n2840), .B(n2841), .C(n2842), .D(n2843), .Y(n2839) );
  AOI22X1 U1846 ( .A0(n18197), .A1(\RAM<55><22> ), .B0(n18189), .B1(
        \RAM<52><22> ), .Y(n2840) );
  AOI22X1 U1847 ( .A0(n18225), .A1(\RAM<53><22> ), .B0(n18218), .B1(
        \RAM<49><22> ), .Y(n2842) );
  AOI22X1 U1848 ( .A0(n18212), .A1(\RAM<51><22> ), .B0(n18204), .B1(
        \RAM<54><22> ), .Y(n2841) );
  NAND4X1 U1849 ( .A(n2860), .B(n2861), .C(n2862), .D(n2863), .Y(n2859) );
  AOI22X1 U1850 ( .A0(n18197), .A1(\RAM<23><22> ), .B0(n18190), .B1(
        \RAM<20><22> ), .Y(n2860) );
  AOI22X1 U1851 ( .A0(n18225), .A1(\RAM<21><22> ), .B0(n18218), .B1(
        \RAM<17><22> ), .Y(n2862) );
  AOI22X1 U1852 ( .A0(n18212), .A1(\RAM<19><22> ), .B0(n18204), .B1(
        \RAM<22><22> ), .Y(n2861) );
  NAND4X1 U1853 ( .A(n2786), .B(n2787), .C(n2788), .D(n2789), .Y(n2785) );
  AOI22X1 U1854 ( .A0(n18198), .A1(\RAM<7><23> ), .B0(n18191), .B1(
        \RAM<4><23> ), .Y(n2786) );
  AOI22X1 U1855 ( .A0(n18226), .A1(\RAM<5><23> ), .B0(n18219), .B1(
        \RAM<1><23> ), .Y(n2788) );
  AOI22X1 U1856 ( .A0(n18213), .A1(\RAM<3><23> ), .B0(n18205), .B1(
        \RAM<6><23> ), .Y(n2787) );
  NAND4X1 U1857 ( .A(n2796), .B(n2797), .C(n2798), .D(n2799), .Y(n2795) );
  AOI22X1 U1858 ( .A0(n18198), .A1(\RAM<55><23> ), .B0(n18191), .B1(
        \RAM<52><23> ), .Y(n2796) );
  AOI22X1 U1859 ( .A0(n18226), .A1(\RAM<53><23> ), .B0(n18219), .B1(
        \RAM<49><23> ), .Y(n2798) );
  AOI22X1 U1860 ( .A0(n18213), .A1(\RAM<51><23> ), .B0(n18205), .B1(
        \RAM<54><23> ), .Y(n2797) );
  NAND4X1 U1861 ( .A(n2816), .B(n2817), .C(n2818), .D(n2819), .Y(n2815) );
  AOI22X1 U1862 ( .A0(n18198), .A1(\RAM<23><23> ), .B0(n18191), .B1(
        \RAM<20><23> ), .Y(n2816) );
  AOI22X1 U1863 ( .A0(n18226), .A1(\RAM<21><23> ), .B0(n18219), .B1(
        \RAM<17><23> ), .Y(n2818) );
  AOI22X1 U1864 ( .A0(n18213), .A1(\RAM<19><23> ), .B0(n18205), .B1(
        \RAM<22><23> ), .Y(n2817) );
  NAND4X1 U1865 ( .A(n2742), .B(n2743), .C(n2744), .D(n2745), .Y(n2741) );
  AOI22X1 U1866 ( .A0(n18198), .A1(\RAM<7><24> ), .B0(n18191), .B1(
        \RAM<4><24> ), .Y(n2742) );
  AOI22X1 U1867 ( .A0(n18226), .A1(\RAM<5><24> ), .B0(n18219), .B1(
        \RAM<1><24> ), .Y(n2744) );
  AOI22X1 U1868 ( .A0(n18213), .A1(\RAM<3><24> ), .B0(n18205), .B1(
        \RAM<6><24> ), .Y(n2743) );
  NAND4X1 U1869 ( .A(n2752), .B(n2753), .C(n2754), .D(n2755), .Y(n2751) );
  AOI22X1 U1870 ( .A0(n18198), .A1(\RAM<55><24> ), .B0(n18191), .B1(
        \RAM<52><24> ), .Y(n2752) );
  AOI22X1 U1871 ( .A0(n18226), .A1(\RAM<53><24> ), .B0(n18219), .B1(
        \RAM<49><24> ), .Y(n2754) );
  AOI22X1 U1872 ( .A0(n18213), .A1(\RAM<51><24> ), .B0(n18205), .B1(
        \RAM<54><24> ), .Y(n2753) );
  NAND4X1 U1873 ( .A(n2772), .B(n2773), .C(n2774), .D(n2775), .Y(n2771) );
  AOI22X1 U1874 ( .A0(n18198), .A1(\RAM<23><24> ), .B0(n18191), .B1(
        \RAM<20><24> ), .Y(n2772) );
  AOI22X1 U1875 ( .A0(n18226), .A1(\RAM<21><24> ), .B0(n18219), .B1(
        \RAM<17><24> ), .Y(n2774) );
  AOI22X1 U1876 ( .A0(n18213), .A1(\RAM<19><24> ), .B0(n18205), .B1(
        \RAM<22><24> ), .Y(n2773) );
  NAND4X1 U1877 ( .A(n2698), .B(n2699), .C(n2700), .D(n2701), .Y(n2697) );
  AOI22X1 U1878 ( .A0(n18198), .A1(\RAM<7><25> ), .B0(n18191), .B1(
        \RAM<4><25> ), .Y(n2698) );
  AOI22X1 U1879 ( .A0(n18226), .A1(\RAM<5><25> ), .B0(n18219), .B1(
        \RAM<1><25> ), .Y(n2700) );
  AOI22X1 U1880 ( .A0(n18213), .A1(\RAM<3><25> ), .B0(n18205), .B1(
        \RAM<6><25> ), .Y(n2699) );
  NAND4X1 U1881 ( .A(n2708), .B(n2709), .C(n2710), .D(n2711), .Y(n2707) );
  AOI22X1 U1882 ( .A0(n18198), .A1(\RAM<55><25> ), .B0(n18191), .B1(
        \RAM<52><25> ), .Y(n2708) );
  AOI22X1 U1883 ( .A0(n18226), .A1(\RAM<53><25> ), .B0(n18219), .B1(
        \RAM<49><25> ), .Y(n2710) );
  AOI22X1 U1884 ( .A0(n18213), .A1(\RAM<51><25> ), .B0(n18205), .B1(
        \RAM<54><25> ), .Y(n2709) );
  NAND4X1 U1885 ( .A(n2728), .B(n2729), .C(n2730), .D(n2731), .Y(n2727) );
  AOI22X1 U1886 ( .A0(n18198), .A1(\RAM<23><25> ), .B0(n18191), .B1(
        \RAM<20><25> ), .Y(n2728) );
  AOI22X1 U1887 ( .A0(n18226), .A1(\RAM<21><25> ), .B0(n18219), .B1(
        \RAM<17><25> ), .Y(n2730) );
  AOI22X1 U1888 ( .A0(n18213), .A1(\RAM<19><25> ), .B0(n18205), .B1(
        \RAM<22><25> ), .Y(n2729) );
  NAND4X1 U1889 ( .A(n2674), .B(n2675), .C(n2676), .D(n2677), .Y(n2673) );
  AOI22X1 U1890 ( .A0(n18199), .A1(\RAM<39><26> ), .B0(n18191), .B1(
        \RAM<36><26> ), .Y(n2674) );
  AOI22X1 U1891 ( .A0(n18227), .A1(\RAM<37><26> ), .B0(n18217), .B1(
        \RAM<33><26> ), .Y(n2676) );
  AOI22X1 U1892 ( .A0(n18214), .A1(\RAM<35><26> ), .B0(n18205), .B1(
        \RAM<38><26> ), .Y(n2675) );
  NAND4X1 U1893 ( .A(n2664), .B(n2665), .C(n2666), .D(n2667), .Y(n2663) );
  AOI22X1 U1894 ( .A0(n18199), .A1(\RAM<55><26> ), .B0(n18191), .B1(
        \RAM<52><26> ), .Y(n2664) );
  AOI22X1 U1895 ( .A0(n18227), .A1(\RAM<53><26> ), .B0(n18216), .B1(
        \RAM<49><26> ), .Y(n2666) );
  AOI22X1 U1896 ( .A0(n18214), .A1(\RAM<51><26> ), .B0(n18205), .B1(
        \RAM<54><26> ), .Y(n2665) );
  NAND4X1 U1897 ( .A(n2684), .B(n2685), .C(n2686), .D(n2687), .Y(n2683) );
  AOI22X1 U1898 ( .A0(n18199), .A1(\RAM<23><26> ), .B0(n18192), .B1(
        \RAM<20><26> ), .Y(n2684) );
  AOI22X1 U1899 ( .A0(n18227), .A1(\RAM<21><26> ), .B0(n18221), .B1(
        \RAM<17><26> ), .Y(n2686) );
  AOI22X1 U1900 ( .A0(n18214), .A1(\RAM<19><26> ), .B0(n18206), .B1(
        \RAM<22><26> ), .Y(n2685) );
  NAND4X1 U1901 ( .A(n2630), .B(n2631), .C(n2632), .D(n2633), .Y(n2629) );
  AOI22X1 U1902 ( .A0(n18199), .A1(\RAM<39><27> ), .B0(n18192), .B1(
        \RAM<36><27> ), .Y(n2630) );
  AOI22X1 U1903 ( .A0(n18227), .A1(\RAM<37><27> ), .B0(n18216), .B1(
        \RAM<33><27> ), .Y(n2632) );
  AOI22X1 U1904 ( .A0(n18214), .A1(\RAM<35><27> ), .B0(n18206), .B1(
        \RAM<38><27> ), .Y(n2631) );
  NAND4X1 U1905 ( .A(n2620), .B(n2621), .C(n2622), .D(n2623), .Y(n2619) );
  AOI22X1 U1906 ( .A0(n18199), .A1(\RAM<55><27> ), .B0(n18191), .B1(
        \RAM<52><27> ), .Y(n2620) );
  AOI22X1 U1907 ( .A0(n18227), .A1(\RAM<53><27> ), .B0(n18221), .B1(
        \RAM<49><27> ), .Y(n2622) );
  AOI22X1 U1908 ( .A0(n18214), .A1(\RAM<51><27> ), .B0(n18205), .B1(
        \RAM<54><27> ), .Y(n2621) );
  NAND4X1 U1909 ( .A(n2640), .B(n2641), .C(n2642), .D(n2643), .Y(n2639) );
  AOI22X1 U1910 ( .A0(n18199), .A1(\RAM<23><27> ), .B0(n18193), .B1(
        \RAM<20><27> ), .Y(n2640) );
  AOI22X1 U1911 ( .A0(n18227), .A1(\RAM<21><27> ), .B0(n18217), .B1(
        \RAM<17><27> ), .Y(n2642) );
  AOI22X1 U1912 ( .A0(n18214), .A1(\RAM<19><27> ), .B0(n18205), .B1(
        \RAM<22><27> ), .Y(n2641) );
  NAND4X1 U1913 ( .A(n2576), .B(n2577), .C(n2578), .D(n2579), .Y(n2575) );
  AOI22X1 U1914 ( .A0(n18199), .A1(\RAM<55><28> ), .B0(n18188), .B1(
        \RAM<52><28> ), .Y(n2576) );
  AOI22X1 U1915 ( .A0(n18227), .A1(\RAM<53><28> ), .B0(n18216), .B1(
        \RAM<49><28> ), .Y(n2578) );
  AOI22X1 U1916 ( .A0(n18214), .A1(\RAM<51><28> ), .B0(n18207), .B1(
        \RAM<54><28> ), .Y(n2577) );
  NAND4X1 U1917 ( .A(n2586), .B(n2587), .C(n2588), .D(n2589), .Y(n2585) );
  AOI22X1 U1918 ( .A0(n18199), .A1(\RAM<39><28> ), .B0(n18188), .B1(
        \RAM<36><28> ), .Y(n2586) );
  AOI22X1 U1919 ( .A0(n18227), .A1(\RAM<37><28> ), .B0(n18217), .B1(
        \RAM<33><28> ), .Y(n2588) );
  AOI22X1 U1920 ( .A0(n18214), .A1(\RAM<35><28> ), .B0(n18207), .B1(
        \RAM<38><28> ), .Y(n2587) );
  NAND4X1 U1921 ( .A(n2596), .B(n2597), .C(n2598), .D(n2599), .Y(n2595) );
  AOI22X1 U1922 ( .A0(n18199), .A1(\RAM<23><28> ), .B0(n18188), .B1(
        \RAM<20><28> ), .Y(n2596) );
  AOI22X1 U1923 ( .A0(n18227), .A1(\RAM<21><28> ), .B0(n18221), .B1(
        \RAM<17><28> ), .Y(n2598) );
  AOI22X1 U1924 ( .A0(n18214), .A1(\RAM<19><28> ), .B0(n18206), .B1(
        \RAM<22><28> ), .Y(n2597) );
  NAND4X1 U1925 ( .A(n2532), .B(n2533), .C(n2534), .D(n2535), .Y(n2531) );
  AOI22X1 U1926 ( .A0(n18198), .A1(\RAM<55><29> ), .B0(n18191), .B1(
        \RAM<52><29> ), .Y(n2532) );
  AOI22X1 U1927 ( .A0(n2069), .A1(\RAM<53><29> ), .B0(n18220), .B1(
        \RAM<49><29> ), .Y(n2534) );
  AOI22X1 U1928 ( .A0(n18213), .A1(\RAM<51><29> ), .B0(n18206), .B1(
        \RAM<54><29> ), .Y(n2533) );
  NAND4X1 U1929 ( .A(n2542), .B(n2543), .C(n2544), .D(n2545), .Y(n2541) );
  AOI22X1 U1930 ( .A0(n18198), .A1(\RAM<39><29> ), .B0(n2074), .B1(
        \RAM<36><29> ), .Y(n2542) );
  AOI22X1 U1931 ( .A0(n18226), .A1(\RAM<37><29> ), .B0(n18220), .B1(
        \RAM<33><29> ), .Y(n2544) );
  AOI22X1 U1932 ( .A0(n18212), .A1(\RAM<35><29> ), .B0(n18206), .B1(
        \RAM<38><29> ), .Y(n2543) );
  NAND4X1 U1933 ( .A(n2552), .B(n2553), .C(n2554), .D(n2555), .Y(n2551) );
  AOI22X1 U1934 ( .A0(n18198), .A1(\RAM<23><29> ), .B0(n2074), .B1(
        \RAM<20><29> ), .Y(n2552) );
  AOI22X1 U1935 ( .A0(n18228), .A1(\RAM<21><29> ), .B0(n18220), .B1(
        \RAM<17><29> ), .Y(n2554) );
  AOI22X1 U1936 ( .A0(n18209), .A1(\RAM<19><29> ), .B0(n18206), .B1(
        \RAM<22><29> ), .Y(n2553) );
  NAND4X1 U1937 ( .A(n2454), .B(n2455), .C(n2456), .D(n2457), .Y(n2453) );
  AOI22X1 U1938 ( .A0(n18197), .A1(\RAM<39><30> ), .B0(n2074), .B1(
        \RAM<36><30> ), .Y(n2454) );
  AOI22X1 U1939 ( .A0(n18226), .A1(\RAM<37><30> ), .B0(n18220), .B1(
        \RAM<33><30> ), .Y(n2456) );
  AOI22X1 U1940 ( .A0(n18212), .A1(\RAM<35><30> ), .B0(n18206), .B1(
        \RAM<38><30> ), .Y(n2455) );
  NAND4X1 U1941 ( .A(n2444), .B(n2445), .C(n2446), .D(n2447), .Y(n2443) );
  AOI22X1 U1942 ( .A0(n18197), .A1(\RAM<55><30> ), .B0(n2074), .B1(
        \RAM<52><30> ), .Y(n2444) );
  AOI22X1 U1943 ( .A0(n18227), .A1(\RAM<53><30> ), .B0(n18220), .B1(
        \RAM<49><30> ), .Y(n2446) );
  AOI22X1 U1944 ( .A0(n18213), .A1(\RAM<51><30> ), .B0(n18206), .B1(
        \RAM<54><30> ), .Y(n2445) );
  NAND4X1 U1945 ( .A(n2464), .B(n2465), .C(n2466), .D(n2467), .Y(n2463) );
  AOI22X1 U1946 ( .A0(n18199), .A1(\RAM<23><30> ), .B0(n18190), .B1(
        \RAM<20><30> ), .Y(n2464) );
  AOI22X1 U1947 ( .A0(n18226), .A1(\RAM<21><30> ), .B0(n18220), .B1(
        \RAM<17><30> ), .Y(n2466) );
  AOI22X1 U1948 ( .A0(n18212), .A1(\RAM<19><30> ), .B0(n18206), .B1(
        \RAM<22><30> ), .Y(n2465) );
  NAND4X1 U1949 ( .A(n2390), .B(n2391), .C(n2392), .D(n2393), .Y(n2389) );
  AOI22X1 U1950 ( .A0(n18200), .A1(\RAM<7><31> ), .B0(n18192), .B1(
        \RAM<4><31> ), .Y(n2390) );
  AOI22X1 U1951 ( .A0(n18224), .A1(\RAM<5><31> ), .B0(n18219), .B1(
        \RAM<1><31> ), .Y(n2392) );
  AOI22X1 U1952 ( .A0(n18213), .A1(\RAM<3><31> ), .B0(n18202), .B1(
        \RAM<6><31> ), .Y(n2391) );
  NAND4X1 U1953 ( .A(n2400), .B(n2401), .C(n2402), .D(n2403), .Y(n2399) );
  AOI22X1 U1954 ( .A0(n18195), .A1(\RAM<55><31> ), .B0(n18192), .B1(
        \RAM<52><31> ), .Y(n2400) );
  AOI22X1 U1955 ( .A0(n18223), .A1(\RAM<53><31> ), .B0(n18219), .B1(
        \RAM<49><31> ), .Y(n2402) );
  AOI22X1 U1956 ( .A0(n18213), .A1(\RAM<51><31> ), .B0(n18202), .B1(
        \RAM<54><31> ), .Y(n2401) );
  NAND4X1 U1957 ( .A(n2420), .B(n2421), .C(n2422), .D(n2423), .Y(n2419) );
  AOI22X1 U1958 ( .A0(n18195), .A1(\RAM<23><31> ), .B0(n18192), .B1(
        \RAM<20><31> ), .Y(n2420) );
  AOI22X1 U1959 ( .A0(n18223), .A1(\RAM<21><31> ), .B0(n18219), .B1(
        \RAM<17><31> ), .Y(n2422) );
  AOI22X1 U1960 ( .A0(n18213), .A1(\RAM<19><31> ), .B0(n18204), .B1(
        \RAM<22><31> ), .Y(n2421) );
  NAND4X1 U1961 ( .A(n3446), .B(n3447), .C(n3448), .D(n3449), .Y(n3445) );
  AOI22X1 U1962 ( .A0(n18195), .A1(\RAM<7><0> ), .B0(n18188), .B1(\RAM<4><0> ), 
        .Y(n3446) );
  AOI22X1 U1963 ( .A0(n18223), .A1(\RAM<5><0> ), .B0(n2070), .B1(\RAM<1><0> ), 
        .Y(n3448) );
  AOI22X1 U1964 ( .A0(n18209), .A1(\RAM<3><0> ), .B0(n2072), .B1(\RAM<6><0> ), 
        .Y(n3447) );
  NAND4X1 U1965 ( .A(n3456), .B(n3457), .C(n3458), .D(n3459), .Y(n3455) );
  AOI22X1 U1966 ( .A0(n18198), .A1(\RAM<55><0> ), .B0(n18188), .B1(
        \RAM<52><0> ), .Y(n3456) );
  AOI22X1 U1967 ( .A0(n18226), .A1(\RAM<53><0> ), .B0(n18220), .B1(
        \RAM<49><0> ), .Y(n3458) );
  AOI22X1 U1968 ( .A0(n18209), .A1(\RAM<51><0> ), .B0(n18205), .B1(
        \RAM<54><0> ), .Y(n3457) );
  NAND4X1 U1969 ( .A(n3476), .B(n3477), .C(n3478), .D(n3479), .Y(n3475) );
  AOI22X1 U1970 ( .A0(n18197), .A1(\RAM<23><0> ), .B0(n18188), .B1(
        \RAM<20><0> ), .Y(n3476) );
  AOI22X1 U1971 ( .A0(n18226), .A1(\RAM<21><0> ), .B0(n18219), .B1(
        \RAM<17><0> ), .Y(n3478) );
  AOI22X1 U1972 ( .A0(n18209), .A1(\RAM<19><0> ), .B0(n18205), .B1(
        \RAM<22><0> ), .Y(n3477) );
  NAND4X1 U1973 ( .A(n2962), .B(n2963), .C(n2964), .D(n2965), .Y(n2961) );
  AOI22X1 U1974 ( .A0(n2073), .A1(\RAM<7><1> ), .B0(n18189), .B1(\RAM<4><1> ), 
        .Y(n2962) );
  AOI22X1 U1975 ( .A0(n18227), .A1(\RAM<5><1> ), .B0(n18216), .B1(\RAM<1><1> ), 
        .Y(n2964) );
  AOI22X1 U1976 ( .A0(n18214), .A1(\RAM<3><1> ), .B0(n18202), .B1(\RAM<6><1> ), 
        .Y(n2963) );
  NAND4X1 U1977 ( .A(n2972), .B(n2973), .C(n2974), .D(n2975), .Y(n2971) );
  AOI22X1 U1978 ( .A0(n2073), .A1(\RAM<55><1> ), .B0(n18190), .B1(\RAM<52><1> ), .Y(n2972) );
  AOI22X1 U1979 ( .A0(n18223), .A1(\RAM<53><1> ), .B0(n18217), .B1(
        \RAM<49><1> ), .Y(n2974) );
  AOI22X1 U1980 ( .A0(n18214), .A1(\RAM<51><1> ), .B0(n18204), .B1(
        \RAM<54><1> ), .Y(n2973) );
  NAND4X1 U1981 ( .A(n2992), .B(n2993), .C(n2994), .D(n2995), .Y(n2991) );
  AOI22X1 U1982 ( .A0(n18196), .A1(\RAM<23><1> ), .B0(n2074), .B1(\RAM<20><1> ), .Y(n2992) );
  AOI22X1 U1983 ( .A0(n18225), .A1(\RAM<21><1> ), .B0(n18216), .B1(
        \RAM<17><1> ), .Y(n2994) );
  AOI22X1 U1984 ( .A0(n18214), .A1(\RAM<19><1> ), .B0(n18203), .B1(
        \RAM<22><1> ), .Y(n2993) );
  NAND4X1 U1985 ( .A(n2126), .B(n2127), .C(n2128), .D(n2129), .Y(n2125) );
  AOI22X1 U1986 ( .A0(n18200), .A1(\RAM<7><8> ), .B0(n18192), .B1(\RAM<4><8> ), 
        .Y(n2126) );
  AOI22X1 U1987 ( .A0(n18227), .A1(\RAM<5><8> ), .B0(n18218), .B1(\RAM<1><8> ), 
        .Y(n2128) );
  AOI22X1 U1988 ( .A0(n18209), .A1(\RAM<3><8> ), .B0(n18207), .B1(\RAM<6><8> ), 
        .Y(n2127) );
  NAND4X1 U1989 ( .A(n2136), .B(n2137), .C(n2138), .D(n2139), .Y(n2135) );
  AOI22X1 U1990 ( .A0(n18200), .A1(\RAM<55><8> ), .B0(n18190), .B1(
        \RAM<52><8> ), .Y(n2136) );
  AOI22X1 U1991 ( .A0(n18228), .A1(\RAM<53><8> ), .B0(n18219), .B1(
        \RAM<49><8> ), .Y(n2138) );
  AOI22X1 U1992 ( .A0(n18209), .A1(\RAM<51><8> ), .B0(n18204), .B1(
        \RAM<54><8> ), .Y(n2137) );
  NAND4X1 U1993 ( .A(n2156), .B(n2157), .C(n2158), .D(n2159), .Y(n2155) );
  AOI22X1 U1994 ( .A0(n18200), .A1(\RAM<23><8> ), .B0(n18192), .B1(
        \RAM<20><8> ), .Y(n2156) );
  AOI22X1 U1995 ( .A0(n18227), .A1(\RAM<21><8> ), .B0(n18218), .B1(
        \RAM<17><8> ), .Y(n2158) );
  AOI22X1 U1996 ( .A0(n18209), .A1(\RAM<19><8> ), .B0(n18207), .B1(
        \RAM<22><8> ), .Y(n2157) );
  NAND4X1 U1997 ( .A(n2063), .B(n2064), .C(n2065), .D(n2066), .Y(n2061) );
  AOI22X1 U1998 ( .A0(n2073), .A1(\RAM<7><9> ), .B0(n18188), .B1(\RAM<4><9> ), 
        .Y(n2063) );
  AOI22X1 U1999 ( .A0(n18225), .A1(\RAM<5><9> ), .B0(n18221), .B1(\RAM<1><9> ), 
        .Y(n2065) );
  AOI22X1 U2000 ( .A0(n2071), .A1(\RAM<3><9> ), .B0(n18207), .B1(\RAM<6><9> ), 
        .Y(n2064) );
  NAND4X1 U2001 ( .A(n2090), .B(n2091), .C(n2092), .D(n2093), .Y(n2088) );
  AOI22X1 U2002 ( .A0(n18198), .A1(\RAM<55><9> ), .B0(n18193), .B1(
        \RAM<52><9> ), .Y(n2090) );
  AOI22X1 U2003 ( .A0(n2069), .A1(\RAM<53><9> ), .B0(n18221), .B1(\RAM<49><9> ), .Y(n2092) );
  AOI22X1 U2004 ( .A0(n18210), .A1(\RAM<51><9> ), .B0(n18206), .B1(
        \RAM<54><9> ), .Y(n2091) );
  NAND4X1 U2005 ( .A(n2112), .B(n2113), .C(n2114), .D(n2115), .Y(n2110) );
  AOI22X1 U2006 ( .A0(n18197), .A1(\RAM<23><9> ), .B0(n18191), .B1(
        \RAM<20><9> ), .Y(n2112) );
  AOI22X1 U2007 ( .A0(n18225), .A1(\RAM<21><9> ), .B0(n18221), .B1(
        \RAM<17><9> ), .Y(n2114) );
  AOI22X1 U2008 ( .A0(n18214), .A1(\RAM<19><9> ), .B0(n18207), .B1(
        \RAM<22><9> ), .Y(n2113) );
endmodule


module top ( clk, reset, .WriteData({\WriteData<31> , \WriteData<30> , 
        \WriteData<29> , \WriteData<28> , \WriteData<27> , \WriteData<26> , 
        \WriteData<25> , \WriteData<24> , \WriteData<23> , \WriteData<22> , 
        \WriteData<21> , \WriteData<20> , \WriteData<19> , \WriteData<18> , 
        \WriteData<17> , \WriteData<16> , \WriteData<15> , \WriteData<14> , 
        \WriteData<13> , \WriteData<12> , \WriteData<11> , \WriteData<10> , 
        \WriteData<9> , \WriteData<8> , \WriteData<7> , \WriteData<6> , 
        \WriteData<5> , \WriteData<4> , \WriteData<3> , \WriteData<2> , 
        \WriteData<1> , \WriteData<0> }), .Adr({\Adr<31> , \Adr<30> , 
        \Adr<29> , \Adr<28> , \Adr<27> , \Adr<26> , \Adr<25> , \Adr<24> , 
        \Adr<23> , \Adr<22> , \Adr<21> , \Adr<20> , \Adr<19> , \Adr<18> , 
        \Adr<17> , \Adr<16> , \Adr<15> , \Adr<14> , \Adr<13> , \Adr<12> , 
        \Adr<11> , \Adr<10> , \Adr<9> , \Adr<8> , \Adr<7> , \Adr<6> , \Adr<5> , 
        \Adr<4> , \Adr<3> , \Adr<2> , \Adr<1> , \Adr<0> }), MemWrite );
  input clk, reset;
  output \WriteData<31> , \WriteData<30> , \WriteData<29> , \WriteData<28> ,
         \WriteData<27> , \WriteData<26> , \WriteData<25> , \WriteData<24> ,
         \WriteData<23> , \WriteData<22> , \WriteData<21> , \WriteData<20> ,
         \WriteData<19> , \WriteData<18> , \WriteData<17> , \WriteData<16> ,
         \WriteData<15> , \WriteData<14> , \WriteData<13> , \WriteData<12> ,
         \WriteData<11> , \WriteData<10> , \WriteData<9> , \WriteData<8> ,
         \WriteData<7> , \WriteData<6> , \WriteData<5> , \WriteData<4> ,
         \WriteData<3> , \WriteData<2> , \WriteData<1> , \WriteData<0> ,
         \Adr<31> , \Adr<30> , \Adr<29> , \Adr<28> , \Adr<27> , \Adr<26> ,
         \Adr<25> , \Adr<24> , \Adr<23> , \Adr<22> , \Adr<21> , \Adr<20> ,
         \Adr<19> , \Adr<18> , \Adr<17> , \Adr<16> , \Adr<15> , \Adr<14> ,
         \Adr<13> , \Adr<12> , \Adr<11> , \Adr<10> , \Adr<9> , \Adr<8> ,
         \Adr<7> , \Adr<6> , \Adr<5> , \Adr<4> , \Adr<3> , \Adr<2> , \Adr<1> ,
         \Adr<0> , MemWrite;
  wire   \ReadData<31> , \ReadData<30> , \ReadData<29> , \ReadData<28> ,
         \ReadData<27> , \ReadData<26> , \ReadData<25> , \ReadData<24> ,
         \ReadData<23> , \ReadData<22> , \ReadData<21> , \ReadData<20> ,
         \ReadData<19> , \ReadData<18> , \ReadData<17> , \ReadData<16> ,
         \ReadData<15> , \ReadData<14> , \ReadData<13> , \ReadData<12> ,
         \ReadData<11> , \ReadData<10> , \ReadData<9> , \ReadData<8> ,
         \ReadData<7> , \ReadData<6> , \ReadData<5> , \ReadData<4> ,
         \ReadData<3> , \ReadData<2> , \ReadData<1> , \ReadData<0> , n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n599, n601,
         n603, n605, n607, n609, n611, n613, n615, n617, n619, n621, n623,
         n625, n627, n629, n631, n633, n635, n637, n639, n641, n643, n645,
         n647, n649, n651, n653, n655, n657, n659, n661;

  arm arm ( .clk(clk), .reset(reset), .MemWrite(MemWrite), .Adr({\Adr<31> , 
        \Adr<30> , \Adr<29> , \Adr<28> , \Adr<27> , \Adr<26> , \Adr<25> , 
        \Adr<24> , \Adr<23> , \Adr<22> , \Adr<21> , \Adr<20> , \Adr<19> , 
        \Adr<18> , \Adr<17> , \Adr<16> , \Adr<15> , \Adr<14> , \Adr<13> , 
        \Adr<12> , \Adr<11> , \Adr<10> , \Adr<9> , \Adr<8> , \Adr<7> , 
        \Adr<6> , \Adr<5> , \Adr<4> , \Adr<3> , \Adr<2> , \Adr<1> , \Adr<0> }), 
        .WriteData({n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, 
        n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, 
        n684, n685, n686, n687, n688, n689, n690, n691, n692, n693}), 
        .ReadData({\ReadData<31> , \ReadData<30> , \ReadData<29> , 
        \ReadData<28> , \ReadData<27> , \ReadData<26> , \ReadData<25> , 
        \ReadData<24> , \ReadData<23> , \ReadData<22> , \ReadData<21> , 
        \ReadData<20> , \ReadData<19> , \ReadData<18> , \ReadData<17> , 
        \ReadData<16> , \ReadData<15> , \ReadData<14> , \ReadData<13> , 
        \ReadData<12> , \ReadData<11> , \ReadData<10> , \ReadData<9> , 
        \ReadData<8> , \ReadData<7> , \ReadData<6> , \ReadData<5> , 
        \ReadData<4> , \ReadData<3> , \ReadData<2> , \ReadData<1> , 
        \ReadData<0> }) );
  mem mem ( .clk(clk), .we(MemWrite), .a({\Adr<31> , \Adr<30> , \Adr<29> , 
        \Adr<28> , \Adr<27> , \Adr<26> , \Adr<25> , \Adr<24> , \Adr<23> , 
        \Adr<22> , \Adr<21> , \Adr<20> , \Adr<19> , \Adr<18> , \Adr<17> , 
        \Adr<16> , \Adr<15> , \Adr<14> , \Adr<13> , \Adr<12> , \Adr<11> , 
        \Adr<10> , \Adr<9> , \Adr<8> , \Adr<7> , \Adr<6> , \Adr<5> , \Adr<4> , 
        \Adr<3> , \Adr<2> , \Adr<1> , \Adr<0> }), .wd({\WriteData<31> , 
        \WriteData<30> , \WriteData<29> , \WriteData<28> , \WriteData<27> , 
        \WriteData<26> , \WriteData<25> , \WriteData<24> , \WriteData<23> , 
        \WriteData<22> , \WriteData<21> , \WriteData<20> , \WriteData<19> , 
        \WriteData<18> , \WriteData<17> , \WriteData<16> , \WriteData<15> , 
        \WriteData<14> , \WriteData<13> , \WriteData<12> , \WriteData<11> , 
        \WriteData<10> , \WriteData<9> , \WriteData<8> , \WriteData<7> , 
        \WriteData<6> , \WriteData<5> , \WriteData<4> , \WriteData<3> , 
        \WriteData<2> , \WriteData<1> , \WriteData<0> }), .rd({\ReadData<31> , 
        \ReadData<30> , \ReadData<29> , \ReadData<28> , \ReadData<27> , 
        \ReadData<26> , \ReadData<25> , \ReadData<24> , \ReadData<23> , 
        \ReadData<22> , \ReadData<21> , \ReadData<20> , \ReadData<19> , 
        \ReadData<18> , \ReadData<17> , \ReadData<16> , \ReadData<15> , 
        \ReadData<14> , \ReadData<13> , \ReadData<12> , \ReadData<11> , 
        \ReadData<10> , \ReadData<9> , \ReadData<8> , \ReadData<7> , 
        \ReadData<6> , \ReadData<5> , \ReadData<4> , \ReadData<3> , 
        \ReadData<2> , \ReadData<1> , \ReadData<0> }) );
  INVX1 U1 ( .A(n599), .Y(\WriteData<0> ) );
  INVX1 U2 ( .A(n693), .Y(n599) );
  INVX1 U3 ( .A(n601), .Y(\WriteData<1> ) );
  INVX1 U4 ( .A(n692), .Y(n601) );
  INVX1 U5 ( .A(n603), .Y(\WriteData<2> ) );
  INVX1 U6 ( .A(n691), .Y(n603) );
  INVX1 U7 ( .A(n605), .Y(\WriteData<3> ) );
  INVX1 U8 ( .A(n690), .Y(n605) );
  INVX1 U9 ( .A(n607), .Y(\WriteData<4> ) );
  INVX1 U10 ( .A(n689), .Y(n607) );
  INVX1 U11 ( .A(n609), .Y(\WriteData<5> ) );
  INVX1 U12 ( .A(n688), .Y(n609) );
  INVX1 U13 ( .A(n611), .Y(\WriteData<6> ) );
  INVX1 U14 ( .A(n687), .Y(n611) );
  INVX1 U15 ( .A(n613), .Y(\WriteData<7> ) );
  INVX1 U16 ( .A(n686), .Y(n613) );
  INVX1 U17 ( .A(n615), .Y(\WriteData<8> ) );
  INVX1 U18 ( .A(n685), .Y(n615) );
  INVX1 U19 ( .A(n617), .Y(\WriteData<9> ) );
  INVX1 U20 ( .A(n684), .Y(n617) );
  INVX1 U21 ( .A(n619), .Y(\WriteData<10> ) );
  INVX1 U22 ( .A(n683), .Y(n619) );
  INVX1 U23 ( .A(n621), .Y(\WriteData<11> ) );
  INVX1 U24 ( .A(n682), .Y(n621) );
  INVX1 U25 ( .A(n623), .Y(\WriteData<12> ) );
  INVX1 U26 ( .A(n681), .Y(n623) );
  INVX1 U27 ( .A(n625), .Y(\WriteData<13> ) );
  INVX1 U28 ( .A(n680), .Y(n625) );
  INVX1 U29 ( .A(n627), .Y(\WriteData<14> ) );
  INVX1 U30 ( .A(n679), .Y(n627) );
  INVX1 U31 ( .A(n629), .Y(\WriteData<15> ) );
  INVX1 U32 ( .A(n678), .Y(n629) );
  INVX1 U33 ( .A(n631), .Y(\WriteData<16> ) );
  INVX1 U34 ( .A(n677), .Y(n631) );
  INVX1 U35 ( .A(n633), .Y(\WriteData<17> ) );
  INVX1 U36 ( .A(n676), .Y(n633) );
  INVX1 U37 ( .A(n635), .Y(\WriteData<18> ) );
  INVX1 U38 ( .A(n675), .Y(n635) );
  INVX1 U39 ( .A(n637), .Y(\WriteData<19> ) );
  INVX1 U40 ( .A(n674), .Y(n637) );
  INVX1 U41 ( .A(n639), .Y(\WriteData<20> ) );
  INVX1 U42 ( .A(n673), .Y(n639) );
  INVX1 U43 ( .A(n641), .Y(\WriteData<21> ) );
  INVX1 U44 ( .A(n672), .Y(n641) );
  INVX1 U45 ( .A(n643), .Y(\WriteData<22> ) );
  INVX1 U46 ( .A(n671), .Y(n643) );
  INVX1 U47 ( .A(n645), .Y(\WriteData<23> ) );
  INVX1 U48 ( .A(n670), .Y(n645) );
  INVX1 U49 ( .A(n647), .Y(\WriteData<24> ) );
  INVX1 U50 ( .A(n669), .Y(n647) );
  INVX1 U51 ( .A(n649), .Y(\WriteData<25> ) );
  INVX1 U52 ( .A(n668), .Y(n649) );
  INVX1 U53 ( .A(n651), .Y(\WriteData<26> ) );
  INVX1 U54 ( .A(n667), .Y(n651) );
  INVX1 U55 ( .A(n653), .Y(\WriteData<27> ) );
  INVX1 U56 ( .A(n666), .Y(n653) );
  INVX1 U57 ( .A(n655), .Y(\WriteData<28> ) );
  INVX1 U58 ( .A(n665), .Y(n655) );
  INVX1 U59 ( .A(n657), .Y(\WriteData<29> ) );
  INVX1 U60 ( .A(n664), .Y(n657) );
  INVX1 U61 ( .A(n659), .Y(\WriteData<30> ) );
  INVX1 U62 ( .A(n663), .Y(n659) );
  INVX1 U63 ( .A(n661), .Y(\WriteData<31> ) );
  INVX1 U64 ( .A(n662), .Y(n661) );
endmodule

